    .INIT_00(256'h022bfc01c002b04f022bfc205062b80f022bfc204fc2b40f022bfc205302b20f),
    .INIT_01(256'h022bfc204d42d010022bfc11c01010e0022bfc14c002b10f022bfc0d5042b08f),
    .INIT_02(256'h022bfc2053e2f032022bfc2054001001022bfc250002d010022bfc204fa0101c),
    .INIT_03(256'h022bfc09c0c204fc022bfc2b03c20500022bfc2b80c20520022bfc204fc2058a),
    .INIT_04(256'h022bfc204d4204fa022bfc09c0c2052e022bfc2b02c20536022bfc204d42200a),
    .INIT_05(256'h022bfc2b00c2051a022bfc204d42051e022bfc09c0c2052a022bfc2b01c25000),
    .INIT_06(256'h022bfc250002052a022bfc204fa25000022bfc204d4204fc022bfc09c0c20538),
    .INIT_07(256'h022bfc20548204fc022bfc2054820540022bfc205482052a022bfc2054820534),
    .INIT_08(256'h022bfc205482051c022bfc2054820520022bfc205482053c022bfc2054825000),
    .INIT_09(256'h022bfc3662c20524022bfc1d00025000022bfc0b032204fc022bfc250002052e),
    .INIT_0A(256'h022bfc204fa0300f022bfc2053c09001022bfc20536204fc022bfc2051e2053e),
    .INIT_0B(256'h022bfc2051a2051a022bfc2053025000022bfc2051e204fa022bfc25000204d3),
    .INIT_0C(256'h022bfc1d00003008022bfc0b03209002022bfc25000204fc022bfc204fa20524),
    .INIT_0D(256'h022bfc20520204d3022bfc205341400e022bfc205221400e022bfc366391400e),
    .INIT_0E(256'h022bfc2051e01100022bfc20522010c0022bfc2500025000022bfc204fa204fa),
    .INIT_0F(256'h022bfc2053801d00022bfc2060a01e02022bfc204fa01f00022bfc2051e207cc),
    .INIT_10(256'h022bfc1410601000022bfc0b11325000022bfc204fc207fa022bfc2051a01c00),
    .INIT_11(256'h022bfc0b00f01e00022bfc1410601f00022bfc14106207cc022bfc1410601103),
    .INIT_12(256'h022bfc204d325000022bfc0b00e207fa022bfc204d301c00022bfc0401001d00),
    .INIT_13(256'h022bfc204d301f00022bfc0b00c207cc022bfc204d301100022bfc0b00d010c0),
    .INIT_14(256'h022bfc204fc207fa022bfc2051a01c00022bfc2053001d01022bfc204fa01e00),
    .INIT_15(256'h022bfc14106207cc022bfc0b11301100022bfc204d3010a0022bfc0100025000),
    .INIT_16(256'h022bfc204d301c00022bfc0401001d00022bfc0b01201e00022bfc1410601f00),
    .INIT_17(256'h022bfc204d303f81022bfc0b010207ea022bfc204d325000022bfc0b011207fa),
    .INIT_18(256'h022bfc1dcff05f00022bfc0bc1703c3f022bfc2500003d7c022bfc204fa03e3c),
    .INIT_19(256'h022bfc346a6207fa022bfc1dcff05c00022bfc0bc1605d02022bfc346a005e40),
    .INIT_1A(256'h022bfc0bc1803e7f022bfc346a003fff022bfc1dcff207ea022bfc0bc1925000),
    .INIT_1B(256'h022bfc1dcff05e80022bfc0bc1b05f00022bfc346a603cff022bfc1dcff03dfd),
    .INIT_1C(256'h022bfc346a625000022bfc1dcff207fa022bfc0bc1a05c00022bfc346a005d00),
    .INIT_1D(256'h022bfc0bc1c25000022bfc346a0207cc022bfc1dcff01101022bfc0bc1d010c0),
    .INIT_1E(256'h022bfc0bd2003dfe022bfc2500003eff022bfc346a603fff022bfc1dcff207ea),
    .INIT_1F(256'h022bfc206a0206b8022bfc0bc1725000022bfc32684207fa022bfc1dd0003cff),
    .INIT_20(256'h022bfc206b220278022bfc0bc2001100022bfc206ac01010022bfc0bc1620274),
    .INIT_21(256'h022bfc0bc1925000022bfc3268d207e3022bfc1dd0001010022bfc0bd2101100),
    .INIT_22(256'h022bfc0bc2101100022bfc206ac01014022bfc0bc1820274022bfc206a0207ae),
    .INIT_23(256'h022bfc32696207e3022bfc1dd0001014022bfc0bd2201100022bfc206b220278),
    .INIT_24(256'h022bfc206ac01018022bfc0bc1a20274022bfc206a0207b4022bfc0bc1b25000),
    .INIT_25(256'h022bfc1dd0001018022bfc0bd2301100022bfc206b220278022bfc0bc2201100),
    .INIT_26(256'h022bfc0bc1c20274022bfc206a0207be022bfc0bc1d25000022bfc3269f207e3),
    .INIT_27(256'h022bfc250000101c022bfc206b220278022bfc0bc2301100022bfc206ac0101c),
    .INIT_28(256'h022bfc204d4207ea022bfc204fc25000022bfc20520207e3022bfc2054601100),
    .INIT_29(256'h022bfc2054003cff022bfc2051c03dfe022bfc2500003eff022bfc204fc03fff),
    .INIT_2A(256'h022bfc2500005c00022bfc204fa05d01022bfc204d405e00022bfc204fc05f00),
    .INIT_2B(256'h022bfc204d420274022bfc204fc206b8022bfc2054025000022bfc2051c207fa),
    .INIT_2C(256'h022bfc2054401100022bfc20530202a3022bfc2500001100022bfc204fc01010),
    .INIT_2D(256'h022bfc25000207ae022bfc204fa25000022bfc204d4207e3022bfc204fc01010),
    .INIT_2E(256'h022bfc2b08e202a3022bfc2b1bb01100022bfc2b21a01014022bfc2bec920274),
    .INIT_2F(256'h022bfc01c0025000022bfc25000207e3022bfc2007301014022bfc2083d01100),
    .INIT_30(256'h022bfc206d101100022bfc01c1001018022bfc2500020274022bfc206d1207b4),
    .INIT_31(256'h022bfc25000207e3022bfc206d101018022bfc01c0701100022bfc25000202a3),
    .INIT_32(256'h022bfc01c010101c022bfc2500020274022bfc206d1207be022bfc01c0d25000),
    .INIT_33(256'h022bfc206d101100022bfc01c040101c022bfc25000202a3022bfc206d101100),
    .INIT_34(256'h022bfc01f001d001022bfc01e000b01e022bfc01d0025000022bfc25000207e3),
    .INIT_35(256'h022bfc207cc0b517022bfc011000b416022bfc0108001200022bfc207d53633b),
    .INIT_36(256'h022bfc2b00a04210022bfc2b3892f917022bfc250002f816022bfc206e020851),
    .INIT_37(256'h022bfc250002f818022bfc2083d20851022bfc2b08e0b519022bfc2b63b0b418),
    .INIT_38(256'h022bfc2b08e0b51b022bfc2b37b0b41a022bfc2b00a04210022bfc2b2092f919),
    .INIT_39(256'h022bfc2b64904210022bfc206ce2f91b022bfc250002f81a022bfc2083d20851),
    .INIT_3A(256'h022bfc2083d2f81c022bfc2b08e20851022bfc2b5bb0b51d022bfc2b62a0b41c),
    .INIT_3B(256'h022bfc206b8322fd022bfc2076e0d202022bfc206b804210022bfc250002f91d),
    .INIT_3C(256'h022bfc2b5bb20625022bfc2b62a2063a022bfc2b6492f21e022bfc206ce01202),
    .INIT_3D(256'h022bfc206b832380022bfc250001d001022bfc2083d0b032022bfc2b08e20632),
    .INIT_3E(256'h022bfc206b805020022bfc2076e20559022bfc206b8323a6022bfc2076e1d002),
    .INIT_3F(256'h022bfc2b5bb208b3022bfc2b62a2f21e022bfc2b64901204022bfc206ce2237c),
    .INIT_40(256'h022bfc206b82f115022bfc250002f014022bfc2083d0b117022bfc2b08e0b016),
    .INIT_41(256'h022bfc206b80b018022bfc2076e3449e022bfc206b81f1ff022bfc2076e1d0ff),
    .INIT_42(256'h022bfc2b6491d0ff022bfc206ce2f115022bfc206b82f014022bfc2076e0b119),
    .INIT_43(256'h022bfc2083d0b11b022bfc2b08e0b01a022bfc2b5bb3449e022bfc2b62a1f1ff),
    .INIT_44(256'h022bfc2b10a1f1ff022bfc2b6491d0ff022bfc206cb2f115022bfc250002f014),
    .INIT_45(256'h022bfc2b6c92f014022bfc2083d0b11d022bfc2b08e0b01c022bfc2bdfb3449e),
    .INIT_46(256'h022bfc2083d3449e022bfc2b08e1f1ff022bfc2bebb1d0ff022bfc2b10a2f115),
    .INIT_47(256'h022bfc207f10b013022bfc01ccc3632f022bfc206b81d000022bfc250000b032),
    .INIT_48(256'h022bfc2b6493232a022bfc206cb1d001022bfc206b832328022bfc207621d000),
    .INIT_49(256'h022bfc2083d3232e022bfc2b08e1d003022bfc2bdfb3232c022bfc2b10a1d002),
    .INIT_4A(256'h022bfc2b08e2232f022bfc2bebb2081c022bfc2b10a2232f022bfc2b6c920812),
    .INIT_4B(256'h022bfc01cd82063a022bfc206b820832022bfc250002232f022bfc2083d20827),
    .INIT_4C(256'h022bfc01ccc0b032022bfc206b820632022bfc2076220662022bfc207f120625),
    .INIT_4D(256'h022bfc206cb323a6022bfc206b81d002022bfc2076232380022bfc207f11d001),
    .INIT_4E(256'h022bfc2b08e1d008022bfc2bdfb2237c022bfc2b10a030df022bfc2b64920559),
    .INIT_4F(256'h022bfc2bebb2051e022bfc2b10a2053c022bfc2b6c92051e022bfc2083d36348),
    .INIT_50(256'h022bfc206b81d001022bfc250000b032022bfc2083d2060a022bfc2b08e204fa),
    .INIT_51(256'h022bfc206b82237c022bfc2076205020022bfc207f120559022bfc01ce432380),
    .INIT_52(256'h022bfc206b820542022bfc207622051a022bfc207f136355022bfc01cd81d010),
    .INIT_53(256'h022bfc206b80b032022bfc207622060a022bfc207f1204fa022bfc01ccc20548),
    .INIT_54(256'h022bfc2bdfb05020022bfc2b10a20559022bfc2b64932380022bfc206cb1d001),
    .INIT_55(256'h022bfc2b10a2051a022bfc2b6c936362022bfc2083d1d020022bfc2b08e2237c),
    .INIT_56(256'h022bfc250002060a022bfc2083d204fa022bfc2b08e20548022bfc2bebb20542),
    .INIT_57(256'h022bfc2b08e20559022bfc2b47b32380022bfc2b22a1d001022bfc2b1c90b032),
    .INIT_58(256'h022bfc2b22a3636f022bfc2b4891d040022bfc250002237c022bfc2083d030df),
    .INIT_59(256'h022bfc25000204fa022bfc2083d20548022bfc2b08e20542022bfc2b57b2051a),
    .INIT_5A(256'h022bfc2b08e32380022bfc2b6bb1d001022bfc2b66a0b032022bfc2b5c92060a),
    .INIT_5B(256'h022bfc2b66a1d080022bfc2b6c92237c022bfc25000030df022bfc2083d20559),
    .INIT_5C(256'h022bfc2500020532022bfc2083d20536022bfc2b08e2053c022bfc2b7bb3602a),
    .INIT_5D(256'h022bfc010801d001022bfc206b80b032022bfc2076e2060a022bfc206b8204fa),
    .INIT_5E(256'h022bfc250002237c022bfc206da030df022bfc207cc20559022bfc0110132380),
    .INIT_5F(256'h022bfc207622200a022bfc207f12056e022bfc01c0e01008022bfc206b820562),
    .INIT_60(256'h022bfc206b81d002022bfc250000b002022bfc206bf20288022bfc206b82027f),
    .INIT_61(256'h022bfc206b81d003022bfc207620b002022bfc207f120291022bfc01c1e3238a),
    .INIT_62(256'h022bfc2076201060022bfc207f120774022bfc01c0e2029a022bfc206bf3238a),
    .INIT_63(256'h022bfc206b82d003022bfc250002f032022bfc206bf01000022bfc206b820562),
    .INIT_64(256'h022bfc206b82b04f022bfc207622b08f022bfc207f12b20f022bfc01c2e2b40f),
    .INIT_65(256'h022bfc207622d010022bfc207f101020022bfc01c1e2d010022bfc206bf01040),
    .INIT_66(256'h022bfc207f12d010022bfc01c0e01004022bfc206bf2d010022bfc206b801008),
    .INIT_67(256'h022bfc250002d010022bfc206bf01080022bfc206b82b10f022bfc207622b80f),
    .INIT_68(256'h022bfc1d0032056e022bfc327a701000022bfc1d0022d010022bfc0b00201010),
    .INIT_69(256'h022bfc2077c2d003022bfc327ab01002022bfc1d0042200a022bfc327a92059c),
    .INIT_6A(256'h022bfc2078f3641a022bfc227ac1d004022bfc207830b01e022bfc227ac2200a),
    .INIT_6B(256'h022bfc01c0e20467022bfc206b8323fe022bfc250000d004022bfc0b00209002),
    .INIT_6C(256'h022bfc25000011b3022bfc206b801e40022bfc2076201f0a022bfc207f12048d),
    .INIT_6D(256'h022bfc207622df0a022bfc207f109d07022bfc01c1a20447022bfc206b80120b),
    .INIT_6E(256'h022bfc20762363bf022bfc207f11ce10022bfc01c0e2dd08022bfc206b82de09),
    .INIT_6F(256'h022bfc01c2611e01022bfc206b8223c2022bfc25000363bf022bfc206b81cf20),
    .INIT_70(256'h022bfc01c1a0b117022bfc206b80b016022bfc20762223b5022bfc207f113f00),
    .INIT_71(256'h022bfc01c0e1f1ff022bfc206b81d0ff022bfc207622f115022bfc207f12f014),
    .INIT_72(256'h022bfc250000d0ff022bfc206b801200022bfc207622044f022bfc207f1323ce),
    .INIT_73(256'h022bfc2d1080b119022bfc2d0080b018022bfc2b4192f220022bfc2b00a14200),
    .INIT_74(256'h022bfc2d1081f1ff022bfc2d0081d0ff022bfc2b2592f115022bfc2b00a2f014),
    .INIT_75(256'h022bfc2dc080d0ff022bfc2b28901200022bfc2b00a2044f022bfc25000323da),
    .INIT_76(256'h022bfc250000b11b022bfc2df080b01a022bfc2de082f221022bfc2dd0814200),
    .INIT_77(256'h022bfc09d081f1ff022bfc09c081d0ff022bfc2b2892f115022bfc2b00a2f014),
    .INIT_78(256'h022bfc2d10a0d0ff022bfc2500001200022bfc09f082044f022bfc09e08323e6),
    .INIT_79(256'h022bfc2de080b11d022bfc2dd080b01c022bfc2dc082f222022bfc2d00914200),
    .INIT_7A(256'h022bfc2d0091d0ff022bfc2d10a2f115022bfc250002f014022bfc2df0801200),
    .INIT_7B(256'h022bfc09f0801200022bfc09e082044f022bfc09d08323f3022bfc09c081f1ff),
    .INIT_7C(256'h022bfc2d10a2062d022bfc011022f223022bfc0105014200022bfc250000d0ff),
    .INIT_7D(256'h022bfc206da0b121022bfc250000b020022bfc2dc0820632022bfc2d0092067b),
    .INIT_7E(256'h022bfc206e00b123022bfc207d504010022bfc250000b122022bfc207dc04010),
    .INIT_7F(256'h022bfc250000504002d00320809205590010ff206b83240102bff02500004010),
    .INITP_00(256'h444744c9f053da51d95f5dc8d9dbcdc15d537e5eefd5e058cac547f964f74e6e),
    .INITP_01(256'hf8e34dfc7ef47cdc6a7e6748c672f0dbe375fffdc4617ef34fd16d7644c6cec8),
    .INITP_02(256'hc960cbf3d679ede674c9ce795871e640d5f6c5e4cb6dd679e8e674f0fbc75871),
    .INITP_03(256'hc1fb42fc477fc555e7c0dd79cbdce9c85bf0c6d5744255e147d9e0c0da71f6d1),
    .INITP_04(256'h77cc684461cffdcd7c4bcc72c2e64d7a4afd51ccf3437d46e1c87bd0cce9c567),
    .INITP_05(256'h7afd5fc067c5e772f453d75e477d725ed0db5567f554d15e58687fda53d46adc),
    .INITP_06(256'h6558e5cf53e661f95c5ad65dea5659fdfa6d74fa6bfaf5e1fd79e974fa69fa77),
    .INITP_07(256'hf0cafbf5d076c8e5416b4d6ee649f5e246fd4f6d51f9e2cdf278e05860ed5363),
    .INITP_08(256'h426159ffc4e6d875db4d62637be7eb754e61e4c6e7edc4f146fe44634a75cfe0),
    .INITP_09(256'h46f4db56fcf66bf269dcf9df7bccf6c07cdc675374d0e94940fd62e3787b40e1),
    .INITP_0A(256'hed427df37941e7457d42d0f07470fc7b4e704770c7fadb6752684af6daffcbe0),
    .INITP_0B(256'he2c9644de37150cccc4ef1427e4a69d5f64de54ce37e6d50f3466562f848e357),
    .INITP_0C(256'he0dfd5f154e5ccc9e9416258d3ecd3e5defc534df7ccef5e5ff546f0dcfcd34a),
    .INITP_0D(256'h64d9e05ce957614cff4de0c1fbd5e9cfe84d78f3e1d6fb53e2745a695170d6ea),
    .INITP_0E(256'h675ad1d8fc416df6495bd4f0615c4cd8ed4069ccfdc0704be95af2c1e342e9d3),
    .INITP_0F(256'he0f8ae4feb477bc0e9f3c95f7c455bfd476c6c4446f47542efe6cfccf2714f67),
