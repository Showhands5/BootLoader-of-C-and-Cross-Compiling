    .INIT_00(256'h0207b42056201f01025000030bf2ff000208092055901f000207ae2240328000),
    .INIT_01(256'h02080919001010010207be0b01f200330250002f03b280000208090b00e2df02),
    .INIT_02(256'h0207cc0b0022df02001100202b701f00001020202ae32077025000364162056e),
    .INIT_03(256'h00bc0c0b0022202a00bd0d202c02202a00be0e324132202a00bf0f1d00228000),
    .INIT_04(256'h001080207742202a0207fd202c92202a025000324132202a0207fa1d0032202a),
    .INIT_05(256'h001100010822202a0010002f01f2202a0207cc224442202a001101010022202a),
    .INIT_06(256'h025000324352202a0207111d0022202a0207fa2200a2202a0207ea205842202a),
    .INIT_07(256'h00110132435280000010801d0102df020207ae3243501f010208001d0082202a),
    .INIT_08(256'h0207ea050401d0040011002055932077001004364271d0010207cc1d0202055c),
    .INIT_09(256'h0208031d0402055f02500022444323a902071d010021d0080207fa20562322d2),
    .INIT_0A(256'h0207cc2056220562001101030bf0106000108020559322d20207b43642e1d004),
    .INIT_0B(256'h0207fa3602a205300207ea1d08020528001100224442056e001008010020109f),
    .INIT_0C(256'h0207be01002200370208062056222bfc025000030bf204fa02072e2055920540),
    .INIT_0D(256'h00100c0b002090020207cc20288250000011012027f20063001080224442004a),
    .INIT_0E(256'h0207430b0020d0010207fa202910b0000207ea3243f320460011001d0020d080),
    .INIT_0F(256'h03683d207740121f00d0082029a011ff00900e3243f010ff0250001d00336046),
    .INIT_10(256'h032841010003e04000d002205621b20000900e050401b1000250002055919001),
    .INIT_11(256'h0328450900d0d04000d0022200a0900100900f2059c2f0000250002056e01001),
    .INIT_12(256'h0328490900d2b00c00d002250002b00000901036447250000250000d08032046),
    .INIT_13(256'h03284d014402d01000d00225000010ff0090113644b2bfff0250000d0402bf7e),
    .INIT_14(256'h00100c0b0142d0010008400b2150300f00095001300090010250000150a2d011),
    .INIT_15(256'h0131000d00809006014808143003605901490e142000d0200011000d0100900d),
    .INIT_16(256'h03685f011010900d01d100030070900603685514300090060190011420022054),
    .INIT_17(256'h00d5082245c2205b02500014106090070018ff3a460360600019ff190010d080),
    .INIT_18(256'h0018ff2d2092053e0019ff2d30a2500000110212350090070368651024009007),
    .INIT_19(256'h00015001a002054203e87225000204fe01d10302010205320250000900820522),
    .INIT_1A(256'h01410e09c1c2051a01180114b062053c0018ff14b06205400000400bb1320530),
    .INIT_1B(256'h00190b10ba0204fe01180809f1f2050403e86a09e1e2054401400809d1d204fe),
    .INIT_1C(256'h00084013f000101900095013e002500002500013d00204fa00110410cb020502),
    .INIT_1D(256'h001102204472022703e87b204912500001b90501b003e07401981801a0419001),
    .INIT_1E(256'h000180204470d00102500009d070900d0018ff20447202150019ff09c072022f),
    .INIT_1F(256'h01410601a730108001490009f07206bf01410620447206b800381f09e073207a),
    .INIT_20(256'h0011020b6121dc930149000b511207f70141060b410207cc01490001b0101101),
    .INIT_21(256'h01400612e60207e301400612d5001000000a9010c4001100000080036013607d),
    .INIT_22(256'h0140063e4851d112014a001bb000311e01400619a01001e001400613f0020898),
    .INIT_23(256'h01d90b204911d11603d00001b01320a201da5d01a741d114014a002500032092),
    .INIT_24(256'h0011042044b2f23903a8952df070122001d8142044b2202a03689325000320b4),
    .INIT_25(256'h0250002044b1400803a8932dd071410a01d8082044b001e00250002de07000d0),
    .INIT_26(256'h0095082044b1d04802f5032db07320c40095082044b1d0580208ac2dc07030f8),
    .INIT_27(256'h009508015001d0b802f6050146c320c702f504250001d0880096082da07320c4),
    .INIT_28(256'h0095080d0102f23902f6310b0140122002f5300b2152202a00960801300320c7),
    .INIT_29(256'h009508142001400802f6380d0081410a02f53714300001e000960814200000d0),
    .INIT_2A(256'h025000190011d08802f60601101320c702f53c030071d04800960814300030f8),
    .INIT_2B(256'h02d509102401d018001100224ab320cc001607141061d0b80015ef3a4af320cc),
    .INIT_2C(256'h001300090082202a0250002d209320ca02d10b2d30a1d00802d60a12350320ca),
    .INIT_2D(256'h02f0162d008001e00208d02d209000d000b1172d30a2f23900b0160601001230),
    .INIT_2E(256'h00b01814c001d08800130114b00030f802f22014a061400802f117250001410a),
    .INIT_2F(256'h02f119250001d0c802f01814f00320c40208d014e001d0b800b11914d00320c4),
    .INIT_30(256'h00b11b14c082202a00b01a14d08320c700130214e081d0e802f22114f0e320c7),
    .INIT_31(256'h02f222110b90100302f11b25000220ce02f01a14a082f0020208d014b0801002),
    .INIT_32(256'h0208d0190112f23900b11d390000124000b01c190e9220ce001303390002f002),
    .INIT_33(256'h025000190f60120302f223390002021102f11d110072f00202f01c3e4d101004),
    .INIT_34(256'h03100000c000100101f1ff250002f03a01d0ff1100a01000001200250002f201),
    .INIT_35(256'h014006204db202550140062054e2024c014006204e520221014006204db2f024),
    .INIT_36(256'h01400e01100207f701410025000202740140062054e20243014100204e52023a),
    .INIT_37(256'h00b224141002027401003014c06207e301400e141000101001400e14c0601100),
    .INIT_38(256'h022bfc1410001100022bfc14c062025e022bfc141000110002500014c0601010),
    .INIT_39(256'h022bfc11107206b8022bfc3a4e8207a0022bfc1d10a207e3022bfc2500001010),
    .INIT_3A(256'h022bfc2055101101022bfc01a0001080022bfc25000206b8022bfc111302076e),
    .INIT_3B(256'h022bfc0110401004022bfc3900001100022bfc204c7207f7022bfc09006207cc),
    .INIT_3C(256'h022bfc04a00207ae022bfc364f02023a022bfc19101207ae022bfc204b9207e3),
    .INIT_3D(256'h022bfc19201207ae022bfc2054e2024c022bfc204e5207ae022bfc0010020243),
    .INIT_3E(256'h022bfc2254e206b8022bfc0110d2076e022bfc25000206b8022bfc364eb20255),
    .INIT_3F(256'h022bfc2254e01014022bfc0115f01100022bfc2254e207f7022bfc0112020274),
    .INIT_40(256'h022bfc2254e207cc022bfc0113101101022bfc2254e010c0022bfc0113e207e3),
    .INIT_41(256'h022bfc2254e2025e022bfc0113001100022bfc2254e01014022bfc01133207ae),
    .INIT_42(256'h022bfc2254e0b002022bfc01132207e3022bfc2254e01014022bfc0113101100),
    .INIT_43(256'h022bfc2254e206b8022bfc01134207a0022bfc2254e32167022bfc011331d002),
    .INIT_44(256'h022bfc2254e206b8022bfc011362076e022bfc2254e206b8022bfc011352076e),
    .INIT_45(256'h022bfc2254e207f7022bfc01138207cc022bfc2254e01101022bfc0113701080),
    .INIT_46(256'h022bfc2254e207b4022bfc01141207e3022bfc2254e01008022bfc0113901100),
    .INIT_47(256'h022bfc2254e207b4022bfc0114320243022bfc2254e207b4022bfc011422023a),
    .INIT_48(256'h022bfc2254e206b8022bfc0114520255022bfc2254e207b4022bfc011442024c),
    .INIT_49(256'h022bfc2254e206b8022bfc011472076e022bfc2254e206b8022bfc011462076e),
    .INIT_4A(256'h022bfc2254e01018022bfc0114901100022bfc2254e207f7022bfc0114820274),
    .INIT_4B(256'h022bfc2254e207cc022bfc0114b01101022bfc2254e010c0022bfc0114a207e3),
    .INIT_4C(256'h022bfc2254e2025e022bfc0114d01100022bfc2254e01018022bfc0114c207b4),
    .INIT_4D(256'h022bfc2254e0b002022bfc0114f207e3022bfc2254e01018022bfc0114e01100),
    .INIT_4E(256'h022bfc2254e206b8022bfc01151207a0022bfc2254e32167022bfc011501d003),
    .INIT_4F(256'h022bfc2254e206b8022bfc011532076e022bfc2254e206b8022bfc011522076e),
    .INIT_50(256'h022bfc2254e01101022bfc0115501080022bfc2254e206b8022bfc011542076e),
    .INIT_51(256'h022bfc2254e0100c022bfc0115701100022bfc2254e207f7022bfc01156207cc),
    .INIT_52(256'h022bfc2254e207be022bfc011592023a022bfc2254e207be022bfc01158207e3),
    .INIT_53(256'h022bfc2d106207be022bfc205552024c022bfc2254e207be022bfc0115a20243),
    .INIT_54(256'h022bfc36551206b8022bfc0d0202076e022bfc0900d206b8022bfc2500020255),
    .INIT_55(256'h022bfc36555206b8022bfc0d0102076e022bfc0900d206b8022bfc250002076e),
    .INIT_56(256'h022bfc250000101c022bfc0306001100022bfc09000207f7022bfc2500020274),
    .INIT_57(256'h022bfc09013207cc022bfc2500001101022bfc0309f010c0022bfc09000207e3),
    .INIT_58(256'h022bfc031602025e022bfc0010001100022bfc250000101c022bfc03007207be),
    .INIT_59(256'h022bfc20524206c5022bfc2d100207e3022bfc041000101c022bfc2055c01100),
    .INIT_5A(256'h022bfc204d3207ae022bfc20559206c5022bfc204fc207ae022bfc2051e206c2),
    .INIT_5B(256'h022bfc0319f3217b022bfc001001d002022bfc250000b002022bfc204fa206c2),
    .INIT_5C(256'h022bfc2053e206c2022bfc2d100207b4022bfc04100206c5022bfc20559207b4),
    .INIT_5D(256'h022bfc1d001207be022bfc0b0323217b022bfc204fc1d003022bfc2051e0b002),
    .INIT_5E(256'h022bfc204fa202ae022bfc204d3206c2022bfc2055c207be022bfc32598206c5),
    .INIT_5F(256'h022bfc204fc32185022bfc2051e1d002022bfc2053e0b002022bfc25000202b7),
    .INIT_60(256'h022bfc2500032185022bfc204fa1d003022bfc204d30b002022bfc01002202c0),
    .INIT_61(256'h022bfc0410001002022bfc205592b02e022bfc0319f20774022bfc00100202c9),
    .INIT_62(256'h022bfc2058401002022bfc010002d010022bfc2500001002022bfc2d1002d00f),
    .INIT_63(256'h022bfc2051e20845022bfc2053e2b02e022bfc2d10320841022bfc0b1322d011),
    .INIT_64(256'h022bfc325981d002022bfc1d0010b002022bfc0b0322d00f022bfc204fc01002),
    .INIT_65(256'h022bfc250002d010022bfc204fa01002022bfc204d320849022bfc010403219e),
    .INIT_66(256'h022bfc250002084d022bfc204fa3219e022bfc204d31d003022bfc010200b002),
    .INIT_67(256'h022bfc205362b02e022bfc325a320841022bfc1d0002d011022bfc2055c01002),
    .INIT_68(256'h022bfc2052a0b002022bfc250002d00f022bfc204fc01002022bfc2050020845),
    .INIT_69(256'h022bfc204fc01002022bfc2053420849022bfc2053e321af022bfc225a01d002),
    .INIT_6A(256'h022bfc20573321af022bfc204fa1d003022bfc204d40b002022bfc00c302d010),
    .INIT_6B(256'h022bfc204fc207a0022bfc2052a2d011022bfc2053c01002022bfc205672084d),
    .INIT_6C(256'h022bfc2500020274022bfc204fa206b8022bfc204d42021b022bfc0bc3a20211),
    .INIT_6D(256'h022bfc2050601100022bfc204fc20269022bfc2052401100022bfc2053201010),
    .INIT_6E(256'h022bfc0bc0520274022bfc204d4207ae022bfc0bc06207e3022bfc2050601010),
    .INIT_6F(256'h022bfc204fa01100022bfc204d420269022bfc0bc0401100022bfc204d401014),
    .INIT_70(256'h022bfc204fc1d002022bfc2051c0b002022bfc20540207e3022bfc2060a01014),
    .INIT_71(256'h022bfc2061c01018022bfc3a5c920274022bfc0d504207b4022bfc09502321d8),
    .INIT_72(256'h022bfc09e1e01018022bfc09d1d01100022bfc09c1c20269022bfc225e001100),
    .INIT_73(256'h022bfc14b06321d8022bfc14b061d003022bfc0bb130b002022bfc09f1f207e3),
    .INIT_74(256'h022bfc13f0001100022bfc13e000101c022bfc13d0020274022bfc10cb0207be),
    .INIT_75(256'h022bfc2fc34207e3022bfc2fd350101c022bfc2fe3601100022bfc2ff3b20269),
    .INIT_76(256'h022bfc204d40300f022bfc0bc3609001022bfc204d42b04e022bfc0bc3b20211),
    .INIT_77(256'h022bfc204d40d002022bfc0bc3409002022bfc204d4321ff022bfc0bc351d001),
    .INIT_78(256'h022bfc204fc2b40f022bfc2051c2b20f022bfc2051e20774022bfc204fa321f0),
    .INIT_79(256'h022bfc225fe2b10f022bfc2061c2b08f022bfc3a5e82b04f022bfc0d5042b80f),
    .INIT_7A(256'h022bfc0bf3b2d010022bfc0be360101c022bfc0bd352d010022bfc0bc34010e0),
    .INIT_7B(256'h022bfc204472200a022bfc204912059c022bfc01b002056e022bfc01a0401002),
    .INIT_7C(256'h022bfc204471d002022bfc09e070b002022bfc2044720288022bfc09f072027f),
    .INIT_7D(256'h022bfc204d41d003022bfc09c070b002022bfc2044720291022bfc09d07321fa),
    .INIT_7E(256'h022bfc204d401000022bfc00ce020774022bfc204d42029a022bfc00cd0321fa),
    .INIT_7F(256'h022bfc2051e20774022bfc204fa2200a022bfc204d42059c022bfc00cf02056e),
    .INITP_00(256'h2c00c765c6f37fda1e09e793b35f5e738ba6a83fd5b53a6d4bdcf84574617be4),
    .INITP_01(256'hce24ac47734bd30784519b8fdde6f57c78f78025691c08d25ac8d6696e842d71),
    .INITP_02(256'h9ce6800dc4a6dc33b20f03b39810afeecfbb1ad04429385bdd0e99585d0b1647),
    .INITP_03(256'hae859fbd2472b9291a5a0eaab0195d2634084e80892223388fc38acd20360073),
    .INITP_04(256'h95f2d6b204738deef6e4bb7b97da87e60a4b31b0aa2ebd27098d112e05b7b70f),
    .INITP_05(256'hfb516311373a4bc0626e840ba8fb68d64f98bf17754ed4b11a45e79e9dddd903),
    .INITP_06(256'h322e8ba8aa0006be9581801057a007bb7e4f6e6f778cb3b3c5c9fb62002233ef),
    .INITP_07(256'heb6b69c3e8ce7372cecd45f8fdf649f2c3dac7585c74737f63f375f6715671da),
    .INITP_08(256'h647f64e96460e35269ca6ac9e853e8d2e84be84b67c1ebcf69d5ebd26b4c6340),
    .INITP_09(256'he8ebe8f1e8f3e8f7677a6aef696e6af96b6a637c6a7269e0e869e873e8726465),
    .INITP_0A(256'hc0f169d27761ddfae8ebc773f46ac7f3f34fe666e66be67965f6696e6aece876),
    .INITP_0B(256'h5361ef7b594e4b53cae646f0eaf6d1cfc9ecfcd643495cf5f2f4df44c2f3774d),
    .INITP_0C(256'heed4cecce25c59e6e0d5d3d7474b7352e973ebddcce5fae75250caf6fbc14b6d),
    .INITP_0D(256'h5d5bea5a78defef97dd9f964fa5cd67d58f27249dac1d6c05271e0f06dee526d),
    .INITP_0E(256'h51f65b68c16bcb67e15251eaf0d6dc547de8c5c8fd78424ee1dfe3c9c56bd479),
    .INITP_0F(256'h74c4565e55c5d948c44d65e6fae968cd7cf1d9617e51c06bdcf542e44ef074d9),
