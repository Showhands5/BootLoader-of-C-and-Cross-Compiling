      parameter integer C_PROBE0_WIDTH         = 1,
      parameter integer C_PROBE1_WIDTH         = 1,
      parameter integer C_PROBE2_WIDTH         = 1,
      parameter integer C_PROBE3_WIDTH         = 1,
      parameter integer C_PROBE4_WIDTH         = 1,
      parameter integer C_PROBE5_WIDTH         = 1,
      parameter integer C_PROBE6_WIDTH         = 1,
      parameter integer C_PROBE7_WIDTH         = 1,
      parameter integer C_PROBE8_WIDTH         = 1,
      parameter integer C_PROBE9_WIDTH         = 1,
      parameter integer C_PROBE10_WIDTH        = 1,
      parameter integer C_PROBE11_WIDTH        = 1,
      parameter integer C_PROBE12_WIDTH        = 1,
      parameter integer C_PROBE13_WIDTH        = 1,
      parameter integer C_PROBE14_WIDTH        = 1,
      parameter integer C_PROBE15_WIDTH        = 1,
      parameter integer C_PROBE16_WIDTH        = 1,
      parameter integer C_PROBE17_WIDTH        = 1,
      parameter integer C_PROBE18_WIDTH        = 1,
      parameter integer C_PROBE19_WIDTH        = 1,
      parameter integer C_PROBE20_WIDTH        = 1,
      parameter integer C_PROBE21_WIDTH        = 1,
      parameter integer C_PROBE22_WIDTH        = 1,
      parameter integer C_PROBE23_WIDTH        = 1,
      parameter integer C_PROBE24_WIDTH        = 1,
      parameter integer C_PROBE25_WIDTH        = 1,
      parameter integer C_PROBE26_WIDTH        = 1,
      parameter integer C_PROBE27_WIDTH        = 1,
      parameter integer C_PROBE28_WIDTH        = 1,
      parameter integer C_PROBE29_WIDTH        = 1,
      parameter integer C_PROBE30_WIDTH        = 1,
      parameter integer C_PROBE31_WIDTH        = 1,
      parameter integer C_PROBE32_WIDTH        = 1,
      parameter integer C_PROBE33_WIDTH        = 1,
      parameter integer C_PROBE34_WIDTH        = 1,
      parameter integer C_PROBE35_WIDTH        = 1,
      parameter integer C_PROBE36_WIDTH        = 1,
      parameter integer C_PROBE37_WIDTH        = 1,
      parameter integer C_PROBE38_WIDTH        = 1,
      parameter integer C_PROBE39_WIDTH        = 1,
      parameter integer C_PROBE40_WIDTH        = 1,
      parameter integer C_PROBE41_WIDTH        = 1,
      parameter integer C_PROBE42_WIDTH        = 1,
      parameter integer C_PROBE43_WIDTH        = 1,
      parameter integer C_PROBE44_WIDTH        = 1,
      parameter integer C_PROBE45_WIDTH        = 1,
      parameter integer C_PROBE46_WIDTH        = 1,
      parameter integer C_PROBE47_WIDTH        = 1,
      parameter integer C_PROBE48_WIDTH        = 1,
      parameter integer C_PROBE49_WIDTH        = 1,
      parameter integer C_PROBE50_WIDTH        = 1,
      parameter integer C_PROBE51_WIDTH        = 1,
      parameter integer C_PROBE52_WIDTH        = 1,
      parameter integer C_PROBE53_WIDTH        = 1,
      parameter integer C_PROBE54_WIDTH        = 1,
      parameter integer C_PROBE55_WIDTH        = 1,
      parameter integer C_PROBE56_WIDTH        = 1,
      parameter integer C_PROBE57_WIDTH        = 1,
      parameter integer C_PROBE58_WIDTH        = 1,
      parameter integer C_PROBE59_WIDTH        = 1,
      parameter integer C_PROBE60_WIDTH        = 1,
      parameter integer C_PROBE61_WIDTH        = 1,
      parameter integer C_PROBE62_WIDTH        = 1,
      parameter integer C_PROBE63_WIDTH        = 1,
      parameter integer C_PROBE64_WIDTH        = 1,
      parameter integer C_PROBE65_WIDTH        = 1,
      parameter integer C_PROBE66_WIDTH        = 1,
      parameter integer C_PROBE67_WIDTH        = 1,
      parameter integer C_PROBE68_WIDTH        = 1,
      parameter integer C_PROBE69_WIDTH        = 1,
      parameter integer C_PROBE70_WIDTH        = 1,
      parameter integer C_PROBE71_WIDTH        = 1,
      parameter integer C_PROBE72_WIDTH        = 1,
      parameter integer C_PROBE73_WIDTH        = 1,
      parameter integer C_PROBE74_WIDTH        = 1,
      parameter integer C_PROBE75_WIDTH        = 1,
      parameter integer C_PROBE76_WIDTH        = 1,
      parameter integer C_PROBE77_WIDTH        = 1,
      parameter integer C_PROBE78_WIDTH        = 1,
      parameter integer C_PROBE79_WIDTH        = 1,
      parameter integer C_PROBE80_WIDTH        = 1,
      parameter integer C_PROBE81_WIDTH        = 1,
      parameter integer C_PROBE82_WIDTH        = 1,
      parameter integer C_PROBE83_WIDTH        = 1,
      parameter integer C_PROBE84_WIDTH        = 1,
      parameter integer C_PROBE85_WIDTH        = 1,
      parameter integer C_PROBE86_WIDTH        = 1,
      parameter integer C_PROBE87_WIDTH        = 1,
      parameter integer C_PROBE88_WIDTH        = 1,
      parameter integer C_PROBE89_WIDTH        = 1,
      parameter integer C_PROBE90_WIDTH        = 1,
      parameter integer C_PROBE91_WIDTH        = 1,
      parameter integer C_PROBE92_WIDTH        = 1,
      parameter integer C_PROBE93_WIDTH        = 1,
      parameter integer C_PROBE94_WIDTH        = 1,
      parameter integer C_PROBE95_WIDTH        = 1,
      parameter integer C_PROBE96_WIDTH        = 1,
      parameter integer C_PROBE97_WIDTH        = 1,
      parameter integer C_PROBE98_WIDTH        = 1,
      parameter integer C_PROBE99_WIDTH        = 1,
      parameter integer C_PROBE100_WIDTH       = 1,
      parameter integer C_PROBE101_WIDTH       = 1,
      parameter integer C_PROBE102_WIDTH       = 1,
      parameter integer C_PROBE103_WIDTH       = 1,
      parameter integer C_PROBE104_WIDTH       = 1,
      parameter integer C_PROBE105_WIDTH       = 1,
      parameter integer C_PROBE106_WIDTH       = 1,
      parameter integer C_PROBE107_WIDTH       = 1,
      parameter integer C_PROBE108_WIDTH       = 1,
      parameter integer C_PROBE109_WIDTH       = 1,
      parameter integer C_PROBE110_WIDTH       = 1,
      parameter integer C_PROBE111_WIDTH       = 1,
      parameter integer C_PROBE112_WIDTH       = 1,
      parameter integer C_PROBE113_WIDTH       = 1,
      parameter integer C_PROBE114_WIDTH       = 1,
      parameter integer C_PROBE115_WIDTH       = 1,
      parameter integer C_PROBE116_WIDTH       = 1,
      parameter integer C_PROBE117_WIDTH       = 1,
      parameter integer C_PROBE118_WIDTH       = 1,
      parameter integer C_PROBE119_WIDTH       = 1,
      parameter integer C_PROBE120_WIDTH       = 1,
      parameter integer C_PROBE121_WIDTH       = 1,
      parameter integer C_PROBE122_WIDTH       = 1,
      parameter integer C_PROBE123_WIDTH       = 1,
      parameter integer C_PROBE124_WIDTH       = 1,
      parameter integer C_PROBE125_WIDTH       = 1,
      parameter integer C_PROBE126_WIDTH       = 1,
      parameter integer C_PROBE127_WIDTH       = 1,
      parameter integer C_PROBE128_WIDTH       = 1,
      parameter integer C_PROBE129_WIDTH       = 1,
      parameter integer C_PROBE130_WIDTH       = 1,
      parameter integer C_PROBE131_WIDTH       = 1,
      parameter integer C_PROBE132_WIDTH       = 1,
      parameter integer C_PROBE133_WIDTH       = 1,
      parameter integer C_PROBE134_WIDTH       = 1,
      parameter integer C_PROBE135_WIDTH       = 1,
      parameter integer C_PROBE136_WIDTH       = 1,
      parameter integer C_PROBE137_WIDTH       = 1,
      parameter integer C_PROBE138_WIDTH       = 1,
      parameter integer C_PROBE139_WIDTH       = 1,
      parameter integer C_PROBE140_WIDTH       = 1,
      parameter integer C_PROBE141_WIDTH       = 1,
      parameter integer C_PROBE142_WIDTH       = 1,
      parameter integer C_PROBE143_WIDTH       = 1,
      parameter integer C_PROBE144_WIDTH       = 1,
      parameter integer C_PROBE145_WIDTH       = 1,
      parameter integer C_PROBE146_WIDTH       = 1,
      parameter integer C_PROBE147_WIDTH       = 1,
      parameter integer C_PROBE148_WIDTH       = 1,
      parameter integer C_PROBE149_WIDTH       = 1,
      parameter integer C_PROBE150_WIDTH       = 1,
      parameter integer C_PROBE151_WIDTH       = 1,
      parameter integer C_PROBE152_WIDTH       = 1,
      parameter integer C_PROBE153_WIDTH       = 1,
      parameter integer C_PROBE154_WIDTH       = 1,
      parameter integer C_PROBE155_WIDTH       = 1,
      parameter integer C_PROBE156_WIDTH       = 1,
      parameter integer C_PROBE157_WIDTH       = 1,
      parameter integer C_PROBE158_WIDTH       = 1,
      parameter integer C_PROBE159_WIDTH       = 1,
      parameter integer C_PROBE160_WIDTH       = 1,
      parameter integer C_PROBE161_WIDTH       = 1,
      parameter integer C_PROBE162_WIDTH       = 1,
      parameter integer C_PROBE163_WIDTH       = 1,
      parameter integer C_PROBE164_WIDTH       = 1,
      parameter integer C_PROBE165_WIDTH       = 1,
      parameter integer C_PROBE166_WIDTH       = 1,
      parameter integer C_PROBE167_WIDTH       = 1,
      parameter integer C_PROBE168_WIDTH       = 1,
      parameter integer C_PROBE169_WIDTH       = 1,
      parameter integer C_PROBE170_WIDTH       = 1,
      parameter integer C_PROBE171_WIDTH       = 1,
      parameter integer C_PROBE172_WIDTH       = 1,
      parameter integer C_PROBE173_WIDTH       = 1,
      parameter integer C_PROBE174_WIDTH       = 1,
      parameter integer C_PROBE175_WIDTH       = 1,
      parameter integer C_PROBE176_WIDTH       = 1,
      parameter integer C_PROBE177_WIDTH       = 1,
      parameter integer C_PROBE178_WIDTH       = 1,
      parameter integer C_PROBE179_WIDTH       = 1,
      parameter integer C_PROBE180_WIDTH       = 1,
      parameter integer C_PROBE181_WIDTH       = 1,
      parameter integer C_PROBE182_WIDTH       = 1,
      parameter integer C_PROBE183_WIDTH       = 1,
      parameter integer C_PROBE184_WIDTH       = 1,
      parameter integer C_PROBE185_WIDTH       = 1,
      parameter integer C_PROBE186_WIDTH       = 1,
      parameter integer C_PROBE187_WIDTH       = 1,
      parameter integer C_PROBE188_WIDTH       = 1,
      parameter integer C_PROBE189_WIDTH       = 1,
      parameter integer C_PROBE190_WIDTH       = 1,
      parameter integer C_PROBE191_WIDTH       = 1,
      parameter integer C_PROBE192_WIDTH       = 1,
      parameter integer C_PROBE193_WIDTH       = 1,
      parameter integer C_PROBE194_WIDTH       = 1,
      parameter integer C_PROBE195_WIDTH       = 1,
      parameter integer C_PROBE196_WIDTH       = 1,
      parameter integer C_PROBE197_WIDTH       = 1,
      parameter integer C_PROBE198_WIDTH       = 1,
      parameter integer C_PROBE199_WIDTH       = 1,
      parameter integer C_PROBE200_WIDTH       = 1,
      parameter integer C_PROBE201_WIDTH       = 1,
      parameter integer C_PROBE202_WIDTH       = 1,
      parameter integer C_PROBE203_WIDTH       = 1,
      parameter integer C_PROBE204_WIDTH       = 1,
      parameter integer C_PROBE205_WIDTH       = 1,
      parameter integer C_PROBE206_WIDTH       = 1,
      parameter integer C_PROBE207_WIDTH       = 1,
      parameter integer C_PROBE208_WIDTH       = 1,
      parameter integer C_PROBE209_WIDTH       = 1,
      parameter integer C_PROBE210_WIDTH       = 1,
      parameter integer C_PROBE211_WIDTH       = 1,
      parameter integer C_PROBE212_WIDTH       = 1,
      parameter integer C_PROBE213_WIDTH       = 1,
      parameter integer C_PROBE214_WIDTH       = 1,
      parameter integer C_PROBE215_WIDTH       = 1,
      parameter integer C_PROBE216_WIDTH       = 1,
      parameter integer C_PROBE217_WIDTH       = 1,
      parameter integer C_PROBE218_WIDTH       = 1,
      parameter integer C_PROBE219_WIDTH       = 1,
      parameter integer C_PROBE220_WIDTH       = 1,
      parameter integer C_PROBE221_WIDTH       = 1,
      parameter integer C_PROBE222_WIDTH       = 1,
      parameter integer C_PROBE223_WIDTH       = 1,
      parameter integer C_PROBE224_WIDTH       = 1,
      parameter integer C_PROBE225_WIDTH       = 1,
      parameter integer C_PROBE226_WIDTH       = 1,
      parameter integer C_PROBE227_WIDTH       = 1,
      parameter integer C_PROBE228_WIDTH       = 1,
      parameter integer C_PROBE229_WIDTH       = 1,
      parameter integer C_PROBE230_WIDTH       = 1,
      parameter integer C_PROBE231_WIDTH       = 1,
      parameter integer C_PROBE232_WIDTH       = 1,
      parameter integer C_PROBE233_WIDTH       = 1,
      parameter integer C_PROBE234_WIDTH       = 1,
      parameter integer C_PROBE235_WIDTH       = 1,
      parameter integer C_PROBE236_WIDTH       = 1,
      parameter integer C_PROBE237_WIDTH       = 1,
      parameter integer C_PROBE238_WIDTH       = 1,
      parameter integer C_PROBE239_WIDTH       = 1,
      parameter integer C_PROBE240_WIDTH       = 1,
      parameter integer C_PROBE241_WIDTH       = 1,
      parameter integer C_PROBE242_WIDTH       = 1,
      parameter integer C_PROBE243_WIDTH       = 1,
      parameter integer C_PROBE244_WIDTH       = 1,
      parameter integer C_PROBE245_WIDTH       = 1,
      parameter integer C_PROBE246_WIDTH       = 1,
      parameter integer C_PROBE247_WIDTH       = 1,
      parameter integer C_PROBE248_WIDTH       = 1,
      parameter integer C_PROBE249_WIDTH       = 1,
      parameter integer C_PROBE250_WIDTH       = 1,
      parameter integer C_PROBE251_WIDTH       = 1,
      parameter integer C_PROBE252_WIDTH       = 1,
      parameter integer C_PROBE253_WIDTH       = 1,
      parameter integer C_PROBE254_WIDTH       = 1,
      parameter integer C_PROBE255_WIDTH       = 1,
