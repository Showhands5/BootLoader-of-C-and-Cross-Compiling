      input  [C_PROBE0_WIDTH-1:0]             probe0,
      input  [C_PROBE1_WIDTH-1:0]             probe1,
      input  [C_PROBE2_WIDTH-1:0]             probe2,
      input  [C_PROBE3_WIDTH-1:0]             probe3,
      input  [C_PROBE4_WIDTH-1:0]             probe4,
      input  [C_PROBE5_WIDTH-1:0]             probe5,
      input  [C_PROBE6_WIDTH-1:0]             probe6,
      input  [C_PROBE7_WIDTH-1:0]             probe7,
      input  [C_PROBE8_WIDTH-1:0]             probe8,
      input  [C_PROBE9_WIDTH-1:0]             probe9,
      input  [C_PROBE10_WIDTH-1:0]            probe10,
      input  [C_PROBE11_WIDTH-1:0]            probe11,
      input  [C_PROBE12_WIDTH-1:0]            probe12,
      input  [C_PROBE13_WIDTH-1:0]            probe13,
      input  [C_PROBE14_WIDTH-1:0]            probe14,
      input  [C_PROBE15_WIDTH-1:0]            probe15,
      input  [C_PROBE16_WIDTH-1:0]            probe16,
      input  [C_PROBE17_WIDTH-1:0]            probe17,
      input  [C_PROBE18_WIDTH-1:0]            probe18,
      input  [C_PROBE19_WIDTH-1:0]            probe19,
      input  [C_PROBE20_WIDTH-1:0]            probe20,
      input  [C_PROBE21_WIDTH-1:0]            probe21,
      input  [C_PROBE22_WIDTH-1:0]            probe22,
      input  [C_PROBE23_WIDTH-1:0]            probe23,
      input  [C_PROBE24_WIDTH-1:0]            probe24,
      input  [C_PROBE25_WIDTH-1:0]            probe25,
      input  [C_PROBE26_WIDTH-1:0]            probe26,
      input  [C_PROBE27_WIDTH-1:0]            probe27,
      input  [C_PROBE28_WIDTH-1:0]            probe28,
      input  [C_PROBE29_WIDTH-1:0]            probe29,
      input  [C_PROBE30_WIDTH-1:0]            probe30,
      input  [C_PROBE31_WIDTH-1:0]            probe31,
      input  [C_PROBE32_WIDTH-1:0]            probe32,
      input  [C_PROBE33_WIDTH-1:0]            probe33,
      input  [C_PROBE34_WIDTH-1:0]            probe34,
      input  [C_PROBE35_WIDTH-1:0]            probe35,
      input  [C_PROBE36_WIDTH-1:0]            probe36,
      input  [C_PROBE37_WIDTH-1:0]            probe37,
      input  [C_PROBE38_WIDTH-1:0]            probe38,
      input  [C_PROBE39_WIDTH-1:0]            probe39,
      input  [C_PROBE40_WIDTH-1:0]            probe40,
      input  [C_PROBE41_WIDTH-1:0]            probe41,
      input  [C_PROBE42_WIDTH-1:0]            probe42,
      input  [C_PROBE43_WIDTH-1:0]            probe43,
      input  [C_PROBE44_WIDTH-1:0]            probe44,
      input  [C_PROBE45_WIDTH-1:0]            probe45,
      input  [C_PROBE46_WIDTH-1:0]            probe46,
      input  [C_PROBE47_WIDTH-1:0]            probe47,
      input  [C_PROBE48_WIDTH-1:0]            probe48,
      input  [C_PROBE49_WIDTH-1:0]            probe49,
      input  [C_PROBE50_WIDTH-1:0]            probe50,
      input  [C_PROBE51_WIDTH-1:0]            probe51,
      input  [C_PROBE52_WIDTH-1:0]            probe52,
      input  [C_PROBE53_WIDTH-1:0]            probe53,
      input  [C_PROBE54_WIDTH-1:0]            probe54,
      input  [C_PROBE55_WIDTH-1:0]            probe55,
      input  [C_PROBE56_WIDTH-1:0]            probe56,
      input  [C_PROBE57_WIDTH-1:0]            probe57,
      input  [C_PROBE58_WIDTH-1:0]            probe58,
      input  [C_PROBE59_WIDTH-1:0]            probe59,
      input  [C_PROBE60_WIDTH-1:0]            probe60,
      input  [C_PROBE61_WIDTH-1:0]            probe61,
      input  [C_PROBE62_WIDTH-1:0]            probe62,
      input  [C_PROBE63_WIDTH-1:0]            probe63,
      input  [C_PROBE64_WIDTH-1:0]            probe64,
      input  [C_PROBE65_WIDTH-1:0]            probe65,
      input  [C_PROBE66_WIDTH-1:0]            probe66,
      input  [C_PROBE67_WIDTH-1:0]            probe67,
      input  [C_PROBE68_WIDTH-1:0]            probe68,
      input  [C_PROBE69_WIDTH-1:0]            probe69,
      input  [C_PROBE70_WIDTH-1:0]            probe70,
      input  [C_PROBE71_WIDTH-1:0]            probe71,
      input  [C_PROBE72_WIDTH-1:0]            probe72,
      input  [C_PROBE73_WIDTH-1:0]            probe73,
      input  [C_PROBE74_WIDTH-1:0]            probe74,
      input  [C_PROBE75_WIDTH-1:0]            probe75,
      input  [C_PROBE76_WIDTH-1:0]            probe76,
      input  [C_PROBE77_WIDTH-1:0]            probe77,
      input  [C_PROBE78_WIDTH-1:0]            probe78,
      input  [C_PROBE79_WIDTH-1:0]            probe79,
      input  [C_PROBE80_WIDTH-1:0]            probe80,
      input  [C_PROBE81_WIDTH-1:0]            probe81,
      input  [C_PROBE82_WIDTH-1:0]            probe82,
      input  [C_PROBE83_WIDTH-1:0]            probe83,
      input  [C_PROBE84_WIDTH-1:0]            probe84,
      input  [C_PROBE85_WIDTH-1:0]            probe85,
      input  [C_PROBE86_WIDTH-1:0]            probe86,
      input  [C_PROBE87_WIDTH-1:0]            probe87,
      input  [C_PROBE88_WIDTH-1:0]            probe88,
      input  [C_PROBE89_WIDTH-1:0]            probe89,
      input  [C_PROBE90_WIDTH-1:0]            probe90,
      input  [C_PROBE91_WIDTH-1:0]            probe91,
      input  [C_PROBE92_WIDTH-1:0]            probe92,
      input  [C_PROBE93_WIDTH-1:0]            probe93,
      input  [C_PROBE94_WIDTH-1:0]            probe94,
      input  [C_PROBE95_WIDTH-1:0]            probe95,
      input  [C_PROBE96_WIDTH-1:0]            probe96,
      input  [C_PROBE97_WIDTH-1:0]            probe97,
      input  [C_PROBE98_WIDTH-1:0]            probe98,
      input  [C_PROBE99_WIDTH-1:0]            probe99,
      input  [C_PROBE100_WIDTH-1:0]           probe100,
      input  [C_PROBE101_WIDTH-1:0]           probe101,
      input  [C_PROBE102_WIDTH-1:0]           probe102,
      input  [C_PROBE103_WIDTH-1:0]           probe103,
      input  [C_PROBE104_WIDTH-1:0]           probe104,
      input  [C_PROBE105_WIDTH-1:0]           probe105,
      input  [C_PROBE106_WIDTH-1:0]           probe106,
      input  [C_PROBE107_WIDTH-1:0]           probe107,
      input  [C_PROBE108_WIDTH-1:0]           probe108,
      input  [C_PROBE109_WIDTH-1:0]           probe109,
      input  [C_PROBE110_WIDTH-1:0]           probe110,
      input  [C_PROBE111_WIDTH-1:0]           probe111,
      input  [C_PROBE112_WIDTH-1:0]           probe112,
      input  [C_PROBE113_WIDTH-1:0]           probe113,
      input  [C_PROBE114_WIDTH-1:0]           probe114,
      input  [C_PROBE115_WIDTH-1:0]           probe115,
      input  [C_PROBE116_WIDTH-1:0]           probe116,
      input  [C_PROBE117_WIDTH-1:0]           probe117,
      input  [C_PROBE118_WIDTH-1:0]           probe118,
      input  [C_PROBE119_WIDTH-1:0]           probe119,
      input  [C_PROBE120_WIDTH-1:0]           probe120,
      input  [C_PROBE121_WIDTH-1:0]           probe121,
      input  [C_PROBE122_WIDTH-1:0]           probe122,
      input  [C_PROBE123_WIDTH-1:0]           probe123,
      input  [C_PROBE124_WIDTH-1:0]           probe124,
      input  [C_PROBE125_WIDTH-1:0]           probe125,
      input  [C_PROBE126_WIDTH-1:0]           probe126,
      input  [C_PROBE127_WIDTH-1:0]           probe127,
      input  [C_PROBE128_WIDTH-1:0]           probe128,
      input  [C_PROBE129_WIDTH-1:0]           probe129,
      input  [C_PROBE130_WIDTH-1:0]           probe130,
      input  [C_PROBE131_WIDTH-1:0]           probe131,
      input  [C_PROBE132_WIDTH-1:0]           probe132,
      input  [C_PROBE133_WIDTH-1:0]           probe133,
      input  [C_PROBE134_WIDTH-1:0]           probe134,
      input  [C_PROBE135_WIDTH-1:0]           probe135,
      input  [C_PROBE136_WIDTH-1:0]           probe136,
      input  [C_PROBE137_WIDTH-1:0]           probe137,
      input  [C_PROBE138_WIDTH-1:0]           probe138,
      input  [C_PROBE139_WIDTH-1:0]           probe139,
      input  [C_PROBE140_WIDTH-1:0]           probe140,
      input  [C_PROBE141_WIDTH-1:0]           probe141,
      input  [C_PROBE142_WIDTH-1:0]           probe142,
      input  [C_PROBE143_WIDTH-1:0]           probe143,
      input  [C_PROBE144_WIDTH-1:0]           probe144,
      input  [C_PROBE145_WIDTH-1:0]           probe145,
      input  [C_PROBE146_WIDTH-1:0]           probe146,
      input  [C_PROBE147_WIDTH-1:0]           probe147,
      input  [C_PROBE148_WIDTH-1:0]           probe148,
      input  [C_PROBE149_WIDTH-1:0]           probe149,
      input  [C_PROBE150_WIDTH-1:0]           probe150,
      input  [C_PROBE151_WIDTH-1:0]           probe151,
      input  [C_PROBE152_WIDTH-1:0]           probe152,
      input  [C_PROBE153_WIDTH-1:0]           probe153,
      input  [C_PROBE154_WIDTH-1:0]           probe154,
      input  [C_PROBE155_WIDTH-1:0]           probe155,
      input  [C_PROBE156_WIDTH-1:0]           probe156,
      input  [C_PROBE157_WIDTH-1:0]           probe157,
      input  [C_PROBE158_WIDTH-1:0]           probe158,
      input  [C_PROBE159_WIDTH-1:0]           probe159,
      input  [C_PROBE160_WIDTH-1:0]           probe160,
      input  [C_PROBE161_WIDTH-1:0]           probe161,
      input  [C_PROBE162_WIDTH-1:0]           probe162,
      input  [C_PROBE163_WIDTH-1:0]           probe163,
      input  [C_PROBE164_WIDTH-1:0]           probe164,
      input  [C_PROBE165_WIDTH-1:0]           probe165,
      input  [C_PROBE166_WIDTH-1:0]           probe166,
      input  [C_PROBE167_WIDTH-1:0]           probe167,
      input  [C_PROBE168_WIDTH-1:0]           probe168,
      input  [C_PROBE169_WIDTH-1:0]           probe169,
      input  [C_PROBE170_WIDTH-1:0]           probe170,
      input  [C_PROBE171_WIDTH-1:0]           probe171,
      input  [C_PROBE172_WIDTH-1:0]           probe172,
      input  [C_PROBE173_WIDTH-1:0]           probe173,
      input  [C_PROBE174_WIDTH-1:0]           probe174,
      input  [C_PROBE175_WIDTH-1:0]           probe175,
      input  [C_PROBE176_WIDTH-1:0]           probe176,
      input  [C_PROBE177_WIDTH-1:0]           probe177,
      input  [C_PROBE178_WIDTH-1:0]           probe178,
      input  [C_PROBE179_WIDTH-1:0]           probe179,
      input  [C_PROBE180_WIDTH-1:0]           probe180,
      input  [C_PROBE181_WIDTH-1:0]           probe181,
      input  [C_PROBE182_WIDTH-1:0]           probe182,
      input  [C_PROBE183_WIDTH-1:0]           probe183,
      input  [C_PROBE184_WIDTH-1:0]           probe184,
      input  [C_PROBE185_WIDTH-1:0]           probe185,
      input  [C_PROBE186_WIDTH-1:0]           probe186,
      input  [C_PROBE187_WIDTH-1:0]           probe187,
      input  [C_PROBE188_WIDTH-1:0]           probe188,
      input  [C_PROBE189_WIDTH-1:0]           probe189,
      input  [C_PROBE190_WIDTH-1:0]           probe190,
      input  [C_PROBE191_WIDTH-1:0]           probe191,
      input  [C_PROBE192_WIDTH-1:0]           probe192,
      input  [C_PROBE193_WIDTH-1:0]           probe193,
      input  [C_PROBE194_WIDTH-1:0]           probe194,
      input  [C_PROBE195_WIDTH-1:0]           probe195,
      input  [C_PROBE196_WIDTH-1:0]           probe196,
      input  [C_PROBE197_WIDTH-1:0]           probe197,
      input  [C_PROBE198_WIDTH-1:0]           probe198,
      input  [C_PROBE199_WIDTH-1:0]           probe199,
      input  [C_PROBE200_WIDTH-1:0]           probe200,
      input  [C_PROBE201_WIDTH-1:0]           probe201,
      input  [C_PROBE202_WIDTH-1:0]           probe202,
      input  [C_PROBE203_WIDTH-1:0]           probe203,
      input  [C_PROBE204_WIDTH-1:0]           probe204,
      input  [C_PROBE205_WIDTH-1:0]           probe205,
      input  [C_PROBE206_WIDTH-1:0]           probe206,
      input  [C_PROBE207_WIDTH-1:0]           probe207,
      input  [C_PROBE208_WIDTH-1:0]           probe208,
      input  [C_PROBE209_WIDTH-1:0]           probe209,
      input  [C_PROBE210_WIDTH-1:0]           probe210,
      input  [C_PROBE211_WIDTH-1:0]           probe211,
      input  [C_PROBE212_WIDTH-1:0]           probe212,
      input  [C_PROBE213_WIDTH-1:0]           probe213,
      input  [C_PROBE214_WIDTH-1:0]           probe214,
      input  [C_PROBE215_WIDTH-1:0]           probe215,
      input  [C_PROBE216_WIDTH-1:0]           probe216,
      input  [C_PROBE217_WIDTH-1:0]           probe217,
      input  [C_PROBE218_WIDTH-1:0]           probe218,
      input  [C_PROBE219_WIDTH-1:0]           probe219,
      input  [C_PROBE220_WIDTH-1:0]           probe220,
      input  [C_PROBE221_WIDTH-1:0]           probe221,
      input  [C_PROBE222_WIDTH-1:0]           probe222,
      input  [C_PROBE223_WIDTH-1:0]           probe223,
      input  [C_PROBE224_WIDTH-1:0]           probe224,
      input  [C_PROBE225_WIDTH-1:0]           probe225,
      input  [C_PROBE226_WIDTH-1:0]           probe226,
      input  [C_PROBE227_WIDTH-1:0]           probe227,
      input  [C_PROBE228_WIDTH-1:0]           probe228,
      input  [C_PROBE229_WIDTH-1:0]           probe229,
      input  [C_PROBE230_WIDTH-1:0]           probe230,
      input  [C_PROBE231_WIDTH-1:0]           probe231,
      input  [C_PROBE232_WIDTH-1:0]           probe232,
      input  [C_PROBE233_WIDTH-1:0]           probe233,
      input  [C_PROBE234_WIDTH-1:0]           probe234,
      input  [C_PROBE235_WIDTH-1:0]           probe235,
      input  [C_PROBE236_WIDTH-1:0]           probe236,
      input  [C_PROBE237_WIDTH-1:0]           probe237,
      input  [C_PROBE238_WIDTH-1:0]           probe238,
      input  [C_PROBE239_WIDTH-1:0]           probe239,
      input  [C_PROBE240_WIDTH-1:0]           probe240,
      input  [C_PROBE241_WIDTH-1:0]           probe241,
      input  [C_PROBE242_WIDTH-1:0]           probe242,
      input  [C_PROBE243_WIDTH-1:0]           probe243,
      input  [C_PROBE244_WIDTH-1:0]           probe244,
      input  [C_PROBE245_WIDTH-1:0]           probe245,
      input  [C_PROBE246_WIDTH-1:0]           probe246,
      input  [C_PROBE247_WIDTH-1:0]           probe247,
      input  [C_PROBE248_WIDTH-1:0]           probe248,
      input  [C_PROBE249_WIDTH-1:0]           probe249,
      input  [C_PROBE250_WIDTH-1:0]           probe250,
      input  [C_PROBE251_WIDTH-1:0]           probe251,
      input  [C_PROBE252_WIDTH-1:0]           probe252,
      input  [C_PROBE253_WIDTH-1:0]           probe253,
      input  [C_PROBE254_WIDTH-1:0]           probe254,
      input  [C_PROBE255_WIDTH-1:0]           probe255,
