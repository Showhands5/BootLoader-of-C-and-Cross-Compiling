   input         cfg_dout0,
   input         cfg_dout1,
   input         cfg_dout2,
   input         cfg_dout3,
   input         cfg_dout4,
   input         cfg_dout5,
   input         cfg_dout6,
   input         cfg_dout7,
   input         cfg_dout8,
   input         cfg_dout9,
   input         cfg_dout10,
   input         cfg_dout11,
   input         cfg_dout12,
   input         cfg_dout13,
   input         cfg_dout14,
   input         cfg_dout15,
   input         cfg_dout16,
   input         cfg_dout17,
   input         cfg_dout18,
   input         cfg_dout19,
   input         cfg_dout20,
   input         cfg_dout21,
   input         cfg_dout22,
   input         cfg_dout23,
   input         cfg_dout24,
   input         cfg_dout25,
   input         cfg_dout26,
   input         cfg_dout27,
   input         cfg_dout28,
   input         cfg_dout29,
   input         cfg_dout30,
   input         cfg_dout31,
   input         cfg_dout32,
   input         cfg_dout33,
   input         cfg_dout34,
   input         cfg_dout35,
   input         cfg_dout36,
   input         cfg_dout37,
   input         cfg_dout38,
   input         cfg_dout39,
   input         cfg_dout40,
   input         cfg_dout41,
   input         cfg_dout42,
   input         cfg_dout43,
   input         cfg_dout44,
   input         cfg_dout45,
   input         cfg_dout46,
   input         cfg_dout47,
   input         cfg_dout48,
   input         cfg_dout49,
   input         cfg_dout50,
   input         cfg_dout51,
   input         cfg_dout52,
   input         cfg_dout53,
   input         cfg_dout54,
   input         cfg_dout55,
   input         cfg_dout56,
   input         cfg_dout57,
   input         cfg_dout58,
   input         cfg_dout59,
   input         cfg_dout60,
   input         cfg_dout61,
   input         cfg_dout62,
   input         cfg_dout63,
   input         cfg_dout64,
   input         cfg_dout65,
   input         cfg_dout66,
   input         cfg_dout67,
   input         cfg_dout68,
   input         cfg_dout69,
   input         cfg_dout70,
   input         cfg_dout71,
   input         cfg_dout72,
   input         cfg_dout73,
   input         cfg_dout74,
   input         cfg_dout75,
   input         cfg_dout76,
   input         cfg_dout77,
   input         cfg_dout78,
   input         cfg_dout79,
   input         cfg_dout80,
   input         cfg_dout81,
   input         cfg_dout82,
   input         cfg_dout83,
   input         cfg_dout84,
   input         cfg_dout85,
   input         cfg_dout86,
   input         cfg_dout87,
   input         cfg_dout88,
   input         cfg_dout89,
   input         cfg_dout90,
   input         cfg_dout91,
   input         cfg_dout92,
   input         cfg_dout93,
   input         cfg_dout94,
   input         cfg_dout95,
   input         cfg_dout96,
   input         cfg_dout97,
   input         cfg_dout98,
   input         cfg_dout99,
   input         cfg_dout100,
   input         cfg_dout101,
   input         cfg_dout102,
   input         cfg_dout103,
   input         cfg_dout104,
   input         cfg_dout105,
   input         cfg_dout106,
   input         cfg_dout107,
   input         cfg_dout108,
   input         cfg_dout109,
   input         cfg_dout110,
   input         cfg_dout111,
   input         cfg_dout112,
   input         cfg_dout113,
   input         cfg_dout114,
   input         cfg_dout115,
   input         cfg_dout116,
   input         cfg_dout117,
   input         cfg_dout118,
   input         cfg_dout119,
   input         cfg_dout120,
   input         cfg_dout121,
   input         cfg_dout122,
   input         cfg_dout123,
   input         cfg_dout124,
   input         cfg_dout125,
   input         cfg_dout126,
   input         cfg_dout127,
   input         cfg_dout128,
   input         cfg_dout129,
   input         cfg_dout130,
   input         cfg_dout131,
   input         cfg_dout132,
   input         cfg_dout133,
   input         cfg_dout134,
   input         cfg_dout135,
   input         cfg_dout136,
   input         cfg_dout137,
   input         cfg_dout138,
   input         cfg_dout139,
   input         cfg_dout140,
   input         cfg_dout141,
   input         cfg_dout142,
   input         cfg_dout143,
   input         cfg_dout144,
   input         cfg_dout145,
   input         cfg_dout146,
   input         cfg_dout147,
   input         cfg_dout148,
   input         cfg_dout149,
   input         cfg_dout150,
   input         cfg_dout151,
   input         cfg_dout152,
   input         cfg_dout153,
   input         cfg_dout154,
   input         cfg_dout155,
   input         cfg_dout156,
   input         cfg_dout157,
   input         cfg_dout158,
   input         cfg_dout159,
   input         cfg_dout160,
   input         cfg_dout161,
   input         cfg_dout162,
   input         cfg_dout163,
   input         cfg_dout164,
   input         cfg_dout165,
   input         cfg_dout166,
   input         cfg_dout167,
   input         cfg_dout168,
   input         cfg_dout169,
   input         cfg_dout170,
   input         cfg_dout171,
   input         cfg_dout172,
   input         cfg_dout173,
   input         cfg_dout174,
   input         cfg_dout175,
   input         cfg_dout176,
   input         cfg_dout177,
   input         cfg_dout178,
   input         cfg_dout179,
   input         cfg_dout180,
   input         cfg_dout181,
   input         cfg_dout182,
   input         cfg_dout183,
   input         cfg_dout184,
   input         cfg_dout185,
   input         cfg_dout186,
   input         cfg_dout187,
   input         cfg_dout188,
   input         cfg_dout189,
   input         cfg_dout190,
   input         cfg_dout191,
   input         cfg_dout192,
   input         cfg_dout193,
   input         cfg_dout194,
   input         cfg_dout195,
   input         cfg_dout196,
   input         cfg_dout197,
   input         cfg_dout198,
   input         cfg_dout199,
   input         cfg_dout200,
   input         cfg_dout201,
   input         cfg_dout202,
   input         cfg_dout203,
   input         cfg_dout204,
   input         cfg_dout205,
   input         cfg_dout206,
   input         cfg_dout207,
   input         cfg_dout208,
   input         cfg_dout209,
   input         cfg_dout210,
   input         cfg_dout211,
   input         cfg_dout212,
   input         cfg_dout213,
   input         cfg_dout214,
   input         cfg_dout215,
   input         cfg_dout216,
   input         cfg_dout217,
   input         cfg_dout218,
   input         cfg_dout219,
   input         cfg_dout220,
   input         cfg_dout221,
   input         cfg_dout222,
   input         cfg_dout223,
   input         cfg_dout224,
   input         cfg_dout225,
   input         cfg_dout226,
   input         cfg_dout227,
   input         cfg_dout228,
   input         cfg_dout229,
   input         cfg_dout230,
   input         cfg_dout231,
   input         cfg_dout232,
   input         cfg_dout233,
   input         cfg_dout234,
   input         cfg_dout235,
   input         cfg_dout236,
   input         cfg_dout237,
   input         cfg_dout238,
   input         cfg_dout239,
   input         cfg_dout240,
   input         cfg_dout241,
   input         cfg_dout242,
   input         cfg_dout243,
   input         cfg_dout244,
   input         cfg_dout245,
   input         cfg_dout246,
   input         cfg_dout247,
   input         cfg_dout248,
   input         cfg_dout249,
   input         cfg_dout250,
   input         cfg_dout251,
   input         cfg_dout252,
   input         cfg_dout253,
   input         cfg_dout254,
   input         cfg_dout255,
   input         cfg_dout256,
   input         cfg_dout257,
   input         cfg_dout258,
   input         cfg_dout259,
   input         cfg_dout260,
   input         cfg_dout261,
   input         cfg_dout262,
   input         cfg_dout263,
   input         cfg_dout264,
   input         cfg_dout265,
   input         cfg_dout266,
   input         cfg_dout267,
   input         cfg_dout268,
   input         cfg_dout269,
   input         cfg_dout270,
   input         cfg_dout271,
   input         cfg_dout272,
   input         cfg_dout273,
   input         cfg_dout274,
   input         cfg_dout275,
   input         cfg_dout276,
   input         cfg_dout277,
   input         cfg_dout278,
   input         cfg_dout279,
   input         cfg_dout280,
   input         cfg_dout281,
   input         cfg_dout282,
   input         cfg_dout283,
   input         cfg_dout284,
   input         cfg_dout285,
   input         cfg_dout286,
   input         cfg_dout287,
   input         cfg_dout288,
   input         cfg_dout289,
   input         cfg_dout290,
   input         cfg_dout291,
   input         cfg_dout292,
   input         cfg_dout293,
   input         cfg_dout294,
   input         cfg_dout295,
   input         cfg_dout296,
   input         cfg_dout297,
   input         cfg_dout298,
   input         cfg_dout299,
   input         cfg_dout300,
   input         cfg_dout301,
   input         cfg_dout302,
   input         cfg_dout303,
   input         cfg_dout304,
   input         cfg_dout305,
   input         cfg_dout306,
   input         cfg_dout307,
   input         cfg_dout308,
   input         cfg_dout309,
   input         cfg_dout310,
   input         cfg_dout311,
   input         cfg_dout312,
   input         cfg_dout313,
   input         cfg_dout314,
   input         cfg_dout315,
   input         cfg_dout316,
   input         cfg_dout317,
   input         cfg_dout318,
   input         cfg_dout319,
   input         cfg_dout320,
   input         cfg_dout321,
   input         cfg_dout322,
   input         cfg_dout323,
   input         cfg_dout324,
   input         cfg_dout325,
   input         cfg_dout326,
   input         cfg_dout327,
   input         cfg_dout328,
   input         cfg_dout329,
   input         cfg_dout330,
   input         cfg_dout331,
   input         cfg_dout332,
   input         cfg_dout333,
   input         cfg_dout334,
   input         cfg_dout335,
   input         cfg_dout336,
   input         cfg_dout337,
   input         cfg_dout338,
   input         cfg_dout339,
   input         cfg_dout340,
   input         cfg_dout341,
   input         cfg_dout342,
   input         cfg_dout343,
   input         cfg_dout344,
   input         cfg_dout345,
   input         cfg_dout346,
   input         cfg_dout347,
   input         cfg_dout348,
   input         cfg_dout349,
   input         cfg_dout350,
   input         cfg_dout351,
   input         cfg_dout352,
   input         cfg_dout353,
   input         cfg_dout354,
   input         cfg_dout355,
   input         cfg_dout356,
   input         cfg_dout357,
   input         cfg_dout358,
   input         cfg_dout359,
   input         cfg_dout360,
   input         cfg_dout361,
   input         cfg_dout362,
   input         cfg_dout363,
   input         cfg_dout364,
   input         cfg_dout365,
   input         cfg_dout366,
   input         cfg_dout367,
   input         cfg_dout368,
   input         cfg_dout369,
   input         cfg_dout370,
   input         cfg_dout371,
   input         cfg_dout372,
   input         cfg_dout373,
   input         cfg_dout374,
   input         cfg_dout375,
   input         cfg_dout376,
   input         cfg_dout377,
   input         cfg_dout378,
   input         cfg_dout379,
   input         cfg_dout380,
   input         cfg_dout381,
   input         cfg_dout382,
   input         cfg_dout383,
   input         cfg_dout384,
   input         cfg_dout385,
   input         cfg_dout386,
   input         cfg_dout387,
   input         cfg_dout388,
   input         cfg_dout389,
   input         cfg_dout390,
   input         cfg_dout391,
   input         cfg_dout392,
   input         cfg_dout393,
   input         cfg_dout394,
   input         cfg_dout395,
   input         cfg_dout396,
   input         cfg_dout397,
   input         cfg_dout398,
   input         cfg_dout399,
   input         cfg_dout400,
   input         cfg_dout401,
   input         cfg_dout402,
   input         cfg_dout403,
   input         cfg_dout404,
   input         cfg_dout405,
   input         cfg_dout406,
   input         cfg_dout407,
   input         cfg_dout408,
   input         cfg_dout409,
   input         cfg_dout410,
   input         cfg_dout411,
   input         cfg_dout412,
   input         cfg_dout413,
   input         cfg_dout414,
   input         cfg_dout415,
   input         cfg_dout416,
   input         cfg_dout417,
   input         cfg_dout418,
   input         cfg_dout419,
   input         cfg_dout420,
   input         cfg_dout421,
   input         cfg_dout422,
   input         cfg_dout423,
   input         cfg_dout424,
   input         cfg_dout425,
   input         cfg_dout426,
   input         cfg_dout427,
   input         cfg_dout428,
   input         cfg_dout429,
   input         cfg_dout430,
   input         cfg_dout431,
   input         cfg_dout432,
   input         cfg_dout433,
   input         cfg_dout434,
   input         cfg_dout435,
   input         cfg_dout436,
   input         cfg_dout437,
   input         cfg_dout438,
   input         cfg_dout439,
   input         cfg_dout440,
   input         cfg_dout441,
   input         cfg_dout442,
   input         cfg_dout443,
   input         cfg_dout444,
   input         cfg_dout445,
   input         cfg_dout446,
   input         cfg_dout447,
   input         cfg_dout448,
   input         cfg_dout449,
   input         cfg_dout450,
   input         cfg_dout451,
   input         cfg_dout452,
   input         cfg_dout453,
   input         cfg_dout454,
   input         cfg_dout455,
   input         cfg_dout456,
   input         cfg_dout457,
   input         cfg_dout458,
   input         cfg_dout459,
   input         cfg_dout460,
   input         cfg_dout461,
   input         cfg_dout462,
   input         cfg_dout463,
   input         cfg_dout464,
   input         cfg_dout465,
   input         cfg_dout466,
   input         cfg_dout467,
   input         cfg_dout468,
   input         cfg_dout469,
   input         cfg_dout470,
   input         cfg_dout471,
   input         cfg_dout472,
   input         cfg_dout473,
   input         cfg_dout474,
   input         cfg_dout475,
   input         cfg_dout476,
   input         cfg_dout477,
   input         cfg_dout478,
   input         cfg_dout479,
   input         cfg_dout480,
   input         cfg_dout481,
   input         cfg_dout482,
   input         cfg_dout483,
   input         cfg_dout484,
   input         cfg_dout485,
   input         cfg_dout486,
   input         cfg_dout487,
   input         cfg_dout488,
   input         cfg_dout489,
   input         cfg_dout490,
   input         cfg_dout491,
   input         cfg_dout492,
   input         cfg_dout493,
   input         cfg_dout494,
   input         cfg_dout495,
   input         cfg_dout496,
   input         cfg_dout497,
   input         cfg_dout498,
   input         cfg_dout499,
   input         cfg_dout500,
   input         cfg_dout501,
   input         cfg_dout502,
   input         cfg_dout503,
   input         cfg_dout504,
   input         cfg_dout505,
   input         cfg_dout506,
   input         cfg_dout507,
   input         cfg_dout508,
   input         cfg_dout509,
   input         cfg_dout510,
   input         cfg_dout511,
   input         cfg_dout512,
   input         cfg_dout513,
   input         cfg_dout514,
   input         cfg_dout515,
   input         cfg_dout516,
   input         cfg_dout517,
   input         cfg_dout518,
   input         cfg_dout519,
   input         cfg_dout520,
   input         cfg_dout521,
   input         cfg_dout522,
   input         cfg_dout523,
   input         cfg_dout524,
   input         cfg_dout525,
   input         cfg_dout526,
   input         cfg_dout527,
   input         cfg_dout528,
   input         cfg_dout529,
   input         cfg_dout530,
   input         cfg_dout531,
   input         cfg_dout532,
   input         cfg_dout533,
   input         cfg_dout534,
   input         cfg_dout535,
   input         cfg_dout536,
   input         cfg_dout537,
   input         cfg_dout538,
   input         cfg_dout539,
   input         cfg_dout540,
   input         cfg_dout541,
   input         cfg_dout542,
   input         cfg_dout543,
   input         cfg_dout544,
   input         cfg_dout545,
   input         cfg_dout546,
   input         cfg_dout547,
   input         cfg_dout548,
   input         cfg_dout549,
   input         cfg_dout550,
   input         cfg_dout551,
   input         cfg_dout552,
   input         cfg_dout553,
   input         cfg_dout554,
   input         cfg_dout555,
   input         cfg_dout556,
   input         cfg_dout557,
   input         cfg_dout558,
   input         cfg_dout559,
   input         cfg_dout560,
   input         cfg_dout561,
   input         cfg_dout562,
   input         cfg_dout563,
   input         cfg_dout564,
   input         cfg_dout565,
   input         cfg_dout566,
   input         cfg_dout567,
   input         cfg_dout568,
   input         cfg_dout569,
   input         cfg_dout570,
   input         cfg_dout571,
   input         cfg_dout572,
   input         cfg_dout573,
   input         cfg_dout574,
   input         cfg_dout575,
   input         cfg_dout576,
   input         cfg_dout577,
   input         cfg_dout578,
   input         cfg_dout579,
   input         cfg_dout580,
   input         cfg_dout581,
   input         cfg_dout582,
   input         cfg_dout583,
   input         cfg_dout584,
   input         cfg_dout585,
   input         cfg_dout586,
   input         cfg_dout587,
   input         cfg_dout588,
   input         cfg_dout589,
   input         cfg_dout590,
   input         cfg_dout591,
   input         cfg_dout592,
   input         cfg_dout593,
   input         cfg_dout594,
   input         cfg_dout595,
   input         cfg_dout596,
   input         cfg_dout597,
   input         cfg_dout598,
   input         cfg_dout599,
   input         cfg_dout600,
   input         cfg_dout601,
   input         cfg_dout602,
   input         cfg_dout603,
   input         cfg_dout604,
   input         cfg_dout605,
   input         cfg_dout606,
   input         cfg_dout607,
   input         cfg_dout608,
   input         cfg_dout609,
   input         cfg_dout610,
   input         cfg_dout611,
   input         cfg_dout612,
   input         cfg_dout613,
   input         cfg_dout614,
   input         cfg_dout615,
   input         cfg_dout616,
   input         cfg_dout617,
   input         cfg_dout618,
   input         cfg_dout619,
   input         cfg_dout620,
   input         cfg_dout621,
   input         cfg_dout622,
   input         cfg_dout623,
   input         cfg_dout624,
   input         cfg_dout625,
   input         cfg_dout626,
   input         cfg_dout627,
   input         cfg_dout628,
   input         cfg_dout629,
   input         cfg_dout630,
   input         cfg_dout631,
   input         cfg_dout632,
   input         cfg_dout633,
   input         cfg_dout634,
   input         cfg_dout635,
   input         cfg_dout636,
   input         cfg_dout637,
   input         cfg_dout638,
   input         cfg_dout639,
   input         cfg_dout640,
   input         cfg_dout641,
   input         cfg_dout642,
   input         cfg_dout643,
   input         cfg_dout644,
   input         cfg_dout645,
   input         cfg_dout646,
   input         cfg_dout647,
   input         cfg_dout648,
   input         cfg_dout649,
   input         cfg_dout650,
   input         cfg_dout651,
   input         cfg_dout652,
   input         cfg_dout653,
   input         cfg_dout654,
   input         cfg_dout655,
   input         cfg_dout656,
   input         cfg_dout657,
   input         cfg_dout658,
   input         cfg_dout659,
   input         cfg_dout660,
   input         cfg_dout661,
   input         cfg_dout662,
   input         cfg_dout663,
   input         cfg_dout664,
   input         cfg_dout665,
   input         cfg_dout666,
   input         cfg_dout667,
   input         cfg_dout668,
   input         cfg_dout669,
   input         cfg_dout670,
   input         cfg_dout671,
   input         cfg_dout672,
   input         cfg_dout673,
   input         cfg_dout674,
   input         cfg_dout675,
   input         cfg_dout676,
   input         cfg_dout677,
   input         cfg_dout678,
   input         cfg_dout679,
   input         cfg_dout680,
   input         cfg_dout681,
   input         cfg_dout682,
   input         cfg_dout683,
   input         cfg_dout684,
   input         cfg_dout685,
   input         cfg_dout686,
   input         cfg_dout687,
   input         cfg_dout688,
   input         cfg_dout689,
   input         cfg_dout690,
   input         cfg_dout691,
   input         cfg_dout692,
   input         cfg_dout693,
   input         cfg_dout694,
   input         cfg_dout695,
   input         cfg_dout696,
   input         cfg_dout697,
   input         cfg_dout698,
   input         cfg_dout699,
   input         cfg_dout700,
   input         cfg_dout701,
   input         cfg_dout702,
   input         cfg_dout703,
   input         cfg_dout704,
   input         cfg_dout705,
   input         cfg_dout706,
   input         cfg_dout707,
   input         cfg_dout708,
   input         cfg_dout709,
   input         cfg_dout710,
   input         cfg_dout711,
   input         cfg_dout712,
   input         cfg_dout713,
   input         cfg_dout714,
   input         cfg_dout715,
   input         cfg_dout716,
   input         cfg_dout717,
   input         cfg_dout718,
   input         cfg_dout719,
   input         cfg_dout720,
   input         cfg_dout721,
   input         cfg_dout722,
   input         cfg_dout723,
   input         cfg_dout724,
   input         cfg_dout725,
   input         cfg_dout726,
   input         cfg_dout727,
   input         cfg_dout728,
   input         cfg_dout729,
   input         cfg_dout730,
   input         cfg_dout731,
   input         cfg_dout732,
   input         cfg_dout733,
   input         cfg_dout734,
   input         cfg_dout735,
   input         cfg_dout736,
   input         cfg_dout737,
   input         cfg_dout738,
   input         cfg_dout739,
   input         cfg_dout740,
   input         cfg_dout741,
   input         cfg_dout742,
   input         cfg_dout743,
   input         cfg_dout744,
   input         cfg_dout745,
   input         cfg_dout746,
   input         cfg_dout747,
   input         cfg_dout748,
   input         cfg_dout749,
   input         cfg_dout750,
   input         cfg_dout751,
   input         cfg_dout752,
   input         cfg_dout753,
   input         cfg_dout754,
   input         cfg_dout755,
   input         cfg_dout756,
   input         cfg_dout757,
   input         cfg_dout758,
   input         cfg_dout759,
   input         cfg_dout760,
   input         cfg_dout761,
   input         cfg_dout762,
   input         cfg_dout763,
   input         cfg_dout764,
   input         cfg_dout765,
   input         cfg_dout766,
   input         cfg_dout767,
   input         cfg_dout768,
   input         cfg_dout769,
   input         cfg_dout770,
   input         cfg_dout771,
   input         cfg_dout772,
   input         cfg_dout773,
   input         cfg_dout774,
   input         cfg_dout775,
   input         cfg_dout776,
   input         cfg_dout777,
   input         cfg_dout778,
   input         cfg_dout779,
   input         cfg_dout780,
   input         cfg_dout781,
   input         cfg_dout782,
   input         cfg_dout783,
   input         cfg_dout784,
   input         cfg_dout785,
   input         cfg_dout786,
   input         cfg_dout787,
   input         cfg_dout788,
   input         cfg_dout789,
   input         cfg_dout790,
   input         cfg_dout791,
   input         cfg_dout792,
   input         cfg_dout793,
   input         cfg_dout794,
   input         cfg_dout795,
   input         cfg_dout796,
   input         cfg_dout797,
   input         cfg_dout798,
   input         cfg_dout799,
   input         cfg_dout800,
   input         cfg_dout801,
   input         cfg_dout802,
   input         cfg_dout803,
   input         cfg_dout804,
   input         cfg_dout805,
   input         cfg_dout806,
   input         cfg_dout807,
   input         cfg_dout808,
   input         cfg_dout809,
   input         cfg_dout810,
   input         cfg_dout811,
   input         cfg_dout812,
   input         cfg_dout813,
   input         cfg_dout814,
   input         cfg_dout815,
   input         cfg_dout816,
   input         cfg_dout817,
   input         cfg_dout818,
   input         cfg_dout819,
   input         cfg_dout820,
   input         cfg_dout821,
   input         cfg_dout822,
   input         cfg_dout823,
   input         cfg_dout824,
   input         cfg_dout825,
   input         cfg_dout826,
   input         cfg_dout827,
   input         cfg_dout828,
   input         cfg_dout829,
   input         cfg_dout830,
   input         cfg_dout831,
   input         cfg_dout832,
   input         cfg_dout833,
   input         cfg_dout834,
   input         cfg_dout835,
   input         cfg_dout836,
   input         cfg_dout837,
   input         cfg_dout838,
   input         cfg_dout839,
   input         cfg_dout840,
   input         cfg_dout841,
   input         cfg_dout842,
   input         cfg_dout843,
   input         cfg_dout844,
   input         cfg_dout845,
   input         cfg_dout846,
   input         cfg_dout847,
   input         cfg_dout848,
   input         cfg_dout849,
   input         cfg_dout850,
   input         cfg_dout851,
   input         cfg_dout852,
   input         cfg_dout853,
   input         cfg_dout854,
   input         cfg_dout855,
   input         cfg_dout856,
   input         cfg_dout857,
   input         cfg_dout858,
   input         cfg_dout859,
   input         cfg_dout860,
   input         cfg_dout861,
   input         cfg_dout862,
   input         cfg_dout863,
   input         cfg_dout864,
   input         cfg_dout865,
   input         cfg_dout866,
   input         cfg_dout867,
   input         cfg_dout868,
   input         cfg_dout869,
   input         cfg_dout870,
   input         cfg_dout871,
   input         cfg_dout872,
   input         cfg_dout873,
   input         cfg_dout874,
   input         cfg_dout875,
   input         cfg_dout876,
   input         cfg_dout877,
   input         cfg_dout878,
   input         cfg_dout879,
   input         cfg_dout880,
   input         cfg_dout881,
   input         cfg_dout882,
   input         cfg_dout883,
   input         cfg_dout884,
   input         cfg_dout885,
   input         cfg_dout886,
   input         cfg_dout887,
   input         cfg_dout888,
   input         cfg_dout889,
   input         cfg_dout890,
   input         cfg_dout891,
   input         cfg_dout892,
   input         cfg_dout893,
   input         cfg_dout894,
   input         cfg_dout895,
   input         cfg_dout896,
   input         cfg_dout897,
   input         cfg_dout898,
   input         cfg_dout899,
   input         cfg_dout900,
   input         cfg_dout901,
   input         cfg_dout902,
   input         cfg_dout903,
   input         cfg_dout904,
   input         cfg_dout905,
   input         cfg_dout906,
   input         cfg_dout907,
   input         cfg_dout908,
   input         cfg_dout909,
   input         cfg_dout910,
   input         cfg_dout911,
   input         cfg_dout912,
   input         cfg_dout913,
   input         cfg_dout914,
   input         cfg_dout915,
   input         cfg_dout916,
   input         cfg_dout917,
   input         cfg_dout918,
   input         cfg_dout919,
   input         cfg_dout920,
   input         cfg_dout921,
   input         cfg_dout922,
   input         cfg_dout923,
   input         cfg_dout924,
   input         cfg_dout925,
   input         cfg_dout926,
   input         cfg_dout927,
   input         cfg_dout928,
   input         cfg_dout929,
   input         cfg_dout930,
   input         cfg_dout931,
   input         cfg_dout932,
   input         cfg_dout933,
   input         cfg_dout934,
   input         cfg_dout935,
   input         cfg_dout936,
   input         cfg_dout937,
   input         cfg_dout938,
   input         cfg_dout939,
   input         cfg_dout940,
   input         cfg_dout941,
   input         cfg_dout942,
   input         cfg_dout943,
   input         cfg_dout944,
   input         cfg_dout945,
   input         cfg_dout946,
   input         cfg_dout947,
   input         cfg_dout948,
   input         cfg_dout949,
   input         cfg_dout950,
   input         cfg_dout951,
   input         cfg_dout952,
   input         cfg_dout953,
   input         cfg_dout954,
   input         cfg_dout955,
   input         cfg_dout956,
   input         cfg_dout957,
   input         cfg_dout958,
   input         cfg_dout959,
   input         cfg_dout960,
   input         cfg_dout961,
   input         cfg_dout962,
   input         cfg_dout963,
   input         cfg_dout964,
   input         cfg_dout965,
   input         cfg_dout966,
   input         cfg_dout967,
   input         cfg_dout968,
   input         cfg_dout969,
   input         cfg_dout970,
   input         cfg_dout971,
   input         cfg_dout972,
   input         cfg_dout973,
   input         cfg_dout974,
   input         cfg_dout975,
   input         cfg_dout976,
   input         cfg_dout977,
   input         cfg_dout978,
   input         cfg_dout979,
   input         cfg_dout980,
   input         cfg_dout981,
   input         cfg_dout982,
   input         cfg_dout983,
   input         cfg_dout984,
   input         cfg_dout985,
   input         cfg_dout986,
   input         cfg_dout987,
   input         cfg_dout988,
   input         cfg_dout989,
   input         cfg_dout990,
   input         cfg_dout991,
   input         cfg_dout992,
   input         cfg_dout993,
   input         cfg_dout994,
   input         cfg_dout995,
   input         cfg_dout996,
   input         cfg_dout997,
   input         cfg_dout998,
   input         cfg_dout999,
   input         cfg_dout1000,
   input         cfg_dout1001,
   input         cfg_dout1002,
   input         cfg_dout1003,
   input         cfg_dout1004,
   input         cfg_dout1005,
   input         cfg_dout1006,
   input         cfg_dout1007,
   input         cfg_dout1008,
   input         cfg_dout1009,
   input         cfg_dout1010,
   input         cfg_dout1011,
   input         cfg_dout1012,
   input         cfg_dout1013,
   input         cfg_dout1014,
   input         cfg_dout1015,
   input         cfg_dout1016,
   input         cfg_dout1017,
   input         cfg_dout1018,
   input         cfg_dout1019,
   input         cfg_dout1020,
   input         cfg_dout1021,
   input         cfg_dout1022,
   input         cfg_dout1023,
   input         cfg_dout1024,
   input         cfg_dout1025,
   input         cfg_dout1026,
   input         cfg_dout1027,
   input         cfg_dout1028,
   input         cfg_dout1029,
   input         cfg_dout1030,
   input         cfg_dout1031,
   input         cfg_dout1032,
   input         cfg_dout1033,
   input         cfg_dout1034,
   input         cfg_dout1035,
   input         cfg_dout1036,
   input         cfg_dout1037,
   input         cfg_dout1038,
   input         cfg_dout1039,
   input         cfg_dout1040,
   input         cfg_dout1041,
   input         cfg_dout1042,
   input         cfg_dout1043,
   input         cfg_dout1044,
   input         cfg_dout1045,
   input         cfg_dout1046,
   input         cfg_dout1047,
   input         cfg_dout1048,
   input         cfg_dout1049,
   input         cfg_dout1050,
   input         cfg_dout1051,
   input         cfg_dout1052,
   input         cfg_dout1053,
   input         cfg_dout1054,
   input         cfg_dout1055,
   input         cfg_dout1056,
   input         cfg_dout1057,
   input         cfg_dout1058,
   input         cfg_dout1059,
   input         cfg_dout1060,
   input         cfg_dout1061,
   input         cfg_dout1062,
   input         cfg_dout1063,
   input         cfg_dout1064,
   input         cfg_dout1065,
   input         cfg_dout1066,
   input         cfg_dout1067,
   input         cfg_dout1068,
   input         cfg_dout1069,
   input         cfg_dout1070,
   input         cfg_dout1071,
   input         cfg_dout1072,
   input         cfg_dout1073,
   input         cfg_dout1074,
   input         cfg_dout1075,
   input         cfg_dout1076,
   input         cfg_dout1077,
   input         cfg_dout1078,
   input         cfg_dout1079,
   input         cfg_dout1080,
   input         cfg_dout1081,
   input         cfg_dout1082,
   input         cfg_dout1083,
   input         cfg_dout1084,
   input         cfg_dout1085,
   input         cfg_dout1086,
   input         cfg_dout1087,
   input         cfg_dout1088,
   input         cfg_dout1089,
   input         cfg_dout1090,
   input         cfg_dout1091,
   input         cfg_dout1092,
   input         cfg_dout1093,
   input         cfg_dout1094,
   input         cfg_dout1095,
   input         cfg_dout1096,
   input         cfg_dout1097,
   input         cfg_dout1098,
   input         cfg_dout1099,
   input         cfg_dout1100,
   input         cfg_dout1101,
   input         cfg_dout1102,
   input         cfg_dout1103,
   input         cfg_dout1104,
   input         cfg_dout1105,
   input         cfg_dout1106,
   input         cfg_dout1107,
   input         cfg_dout1108,
   input         cfg_dout1109,
   input         cfg_dout1110,
   input         cfg_dout1111,
   input         cfg_dout1112,
   input         cfg_dout1113,
   input         cfg_dout1114,
   input         cfg_dout1115,
   input         cfg_dout1116,
   input         cfg_dout1117,
   input         cfg_dout1118,
   input         cfg_dout1119,
   input         cfg_dout1120,
   input         cfg_dout1121,
   input         cfg_dout1122,
   input         cfg_dout1123,
   input         cfg_dout1124,
   input         cfg_dout1125,
   input         cfg_dout1126,
   input         cfg_dout1127,
   input         cfg_dout1128,
   input         cfg_dout1129,
   input         cfg_dout1130,
   input         cfg_dout1131,
   input         cfg_dout1132,
   input         cfg_dout1133,
   input         cfg_dout1134,
   input         cfg_dout1135,
   input         cfg_dout1136,
   input         cfg_dout1137,
   input         cfg_dout1138,
   input         cfg_dout1139,
   input         cfg_dout1140,
   input         cfg_dout1141,
   input         cfg_dout1142,
   input         cfg_dout1143,
   input         cfg_dout1144,
   input         cfg_dout1145,
   input         cfg_dout1146,
   input         cfg_dout1147,
   input         cfg_dout1148,
   input         cfg_dout1149,
   input         cfg_dout1150,
   input         cfg_dout1151,
   input         cfg_dout1152,
   input         cfg_dout1153,
   input         cfg_dout1154,
   input         cfg_dout1155,
   input         cfg_dout1156,
   input         cfg_dout1157,
   input         cfg_dout1158,
   input         cfg_dout1159,
   input         cfg_dout1160,
   input         cfg_dout1161,
   input         cfg_dout1162,
   input         cfg_dout1163,
   input         cfg_dout1164,
   input         cfg_dout1165,
   input         cfg_dout1166,
   input         cfg_dout1167,
   input         cfg_dout1168,
   input         cfg_dout1169,
   input         cfg_dout1170,
   input         cfg_dout1171,
   input         cfg_dout1172,
   input         cfg_dout1173,
   input         cfg_dout1174,
   input         cfg_dout1175,
   input         cfg_dout1176,
   input         cfg_dout1177,
   input         cfg_dout1178,
   input         cfg_dout1179,
   input         cfg_dout1180,
   input         cfg_dout1181,
   input         cfg_dout1182,
   input         cfg_dout1183,
   input         cfg_dout1184,
   input         cfg_dout1185,
   input         cfg_dout1186,
   input         cfg_dout1187,
   input         cfg_dout1188,
   input         cfg_dout1189,
   input         cfg_dout1190,
   input         cfg_dout1191,
   input         cfg_dout1192,
   input         cfg_dout1193,
   input         cfg_dout1194,
   input         cfg_dout1195,
   input         cfg_dout1196,
   input         cfg_dout1197,
   input         cfg_dout1198,
   input         cfg_dout1199,
   input         cfg_dout1200,
   input         cfg_dout1201,
   input         cfg_dout1202,
   input         cfg_dout1203,
   input         cfg_dout1204,
   input         cfg_dout1205,
   input         cfg_dout1206,
   input         cfg_dout1207,
   input         cfg_dout1208,
   input         cfg_dout1209,
   input         cfg_dout1210,
   input         cfg_dout1211,
   input         cfg_dout1212,
   input         cfg_dout1213,
   input         cfg_dout1214,
   input         cfg_dout1215,
   input         cfg_dout1216,
   input         cfg_dout1217,
   input         cfg_dout1218,
   input         cfg_dout1219,
   input         cfg_dout1220,
   input         cfg_dout1221,
   input         cfg_dout1222,
   input         cfg_dout1223,
   input         cfg_dout1224,
   input         cfg_dout1225,
   input         cfg_dout1226,
   input         cfg_dout1227,
   input         cfg_dout1228,
   input         cfg_dout1229,
   input         cfg_dout1230,
   input         cfg_dout1231,
   input         cfg_dout1232,
   input         cfg_dout1233,
   input         cfg_dout1234,
   input         cfg_dout1235,
   input         cfg_dout1236,
   input         cfg_dout1237,
   input         cfg_dout1238,
   input         cfg_dout1239,
   input         cfg_dout1240,
   input         cfg_dout1241,
   input         cfg_dout1242,
   input         cfg_dout1243,
   input         cfg_dout1244,
   input         cfg_dout1245,
   input         cfg_dout1246,
   input         cfg_dout1247,
   input         cfg_dout1248,
   input         cfg_dout1249,
   input         cfg_dout1250,
   input         cfg_dout1251,
   input         cfg_dout1252,
   input         cfg_dout1253,
   input         cfg_dout1254,
   input         cfg_dout1255,
   input         cfg_dout1256,
   input         cfg_dout1257,
   input         cfg_dout1258,
   input         cfg_dout1259,
   input         cfg_dout1260,
   input         cfg_dout1261,
   input         cfg_dout1262,
   input         cfg_dout1263,
   input         cfg_dout1264,
   input         cfg_dout1265,
   input         cfg_dout1266,
   input         cfg_dout1267,
   input         cfg_dout1268,
   input         cfg_dout1269,
   input         cfg_dout1270,
   input         cfg_dout1271,
   input         cfg_dout1272,
   input         cfg_dout1273,
   input         cfg_dout1274,
   input         cfg_dout1275,
   input         cfg_dout1276,
   input         cfg_dout1277,
   input         cfg_dout1278,
   input         cfg_dout1279,
   input         cfg_dout1280,
   input         cfg_dout1281,
   input         cfg_dout1282,
   input         cfg_dout1283,
   input         cfg_dout1284,
   input         cfg_dout1285,
   input         cfg_dout1286,
   input         cfg_dout1287,
   input         cfg_dout1288,
   input         cfg_dout1289,
   input         cfg_dout1290,
   input         cfg_dout1291,
   input         cfg_dout1292,
   input         cfg_dout1293,
   input         cfg_dout1294,
   input         cfg_dout1295,
   input         cfg_dout1296,
   input         cfg_dout1297,
   input         cfg_dout1298,
   input         cfg_dout1299,
   input         cfg_dout1300,
   input         cfg_dout1301,
   input         cfg_dout1302,
   input         cfg_dout1303,
   input         cfg_dout1304,
   input         cfg_dout1305,
   input         cfg_dout1306,
   input         cfg_dout1307,
   input         cfg_dout1308,
   input         cfg_dout1309,
   input         cfg_dout1310,
   input         cfg_dout1311,
   input         cfg_dout1312,
   input         cfg_dout1313,
   input         cfg_dout1314,
   input         cfg_dout1315,
   input         cfg_dout1316,
   input         cfg_dout1317,
   input         cfg_dout1318,
   input         cfg_dout1319,
   input         cfg_dout1320,
   input         cfg_dout1321,
   input         cfg_dout1322,
   input         cfg_dout1323,
   input         cfg_dout1324,
   input         cfg_dout1325,
   input         cfg_dout1326,
   input         cfg_dout1327,
   input         cfg_dout1328,
   input         cfg_dout1329,
   input         cfg_dout1330,
   input         cfg_dout1331,
   input         cfg_dout1332,
   input         cfg_dout1333,
   input         cfg_dout1334,
   input         cfg_dout1335,
   input         cfg_dout1336,
   input         cfg_dout1337,
   input         cfg_dout1338,
   input         cfg_dout1339,
   input         cfg_dout1340,
   input         cfg_dout1341,
   input         cfg_dout1342,
   input         cfg_dout1343,
   input         cfg_dout1344,
   input         cfg_dout1345,
   input         cfg_dout1346,
   input         cfg_dout1347,
   input         cfg_dout1348,
   input         cfg_dout1349,
   input         cfg_dout1350,
   input         cfg_dout1351,
   input         cfg_dout1352,
   input         cfg_dout1353,
   input         cfg_dout1354,
   input         cfg_dout1355,
   input         cfg_dout1356,
   input         cfg_dout1357,
   input         cfg_dout1358,
   input         cfg_dout1359,
   input         cfg_dout1360,
   input         cfg_dout1361,
   input         cfg_dout1362,
   input         cfg_dout1363,
   input         cfg_dout1364,
   input         cfg_dout1365,
   input         cfg_dout1366,
   input         cfg_dout1367,
   input         cfg_dout1368,
   input         cfg_dout1369,
   input         cfg_dout1370,
   input         cfg_dout1371,
   input         cfg_dout1372,
   input         cfg_dout1373,
   input         cfg_dout1374,
   input         cfg_dout1375,
   input         cfg_dout1376,
   input         cfg_dout1377,
   input         cfg_dout1378,
   input         cfg_dout1379,
   input         cfg_dout1380,
   input         cfg_dout1381,
   input         cfg_dout1382,
   input         cfg_dout1383,
   input         cfg_dout1384,
   input         cfg_dout1385,
   input         cfg_dout1386,
   input         cfg_dout1387,
   input         cfg_dout1388,
   input         cfg_dout1389,
   input         cfg_dout1390,
   input         cfg_dout1391,
   input         cfg_dout1392,
   input         cfg_dout1393,
   input         cfg_dout1394,
   input         cfg_dout1395,
   input         cfg_dout1396,
   input         cfg_dout1397,
   input         cfg_dout1398,
   input         cfg_dout1399,
   input         cfg_dout1400,
   input         cfg_dout1401,
   input         cfg_dout1402,
   input         cfg_dout1403,
   input         cfg_dout1404,
   input         cfg_dout1405,
   input         cfg_dout1406,
   input         cfg_dout1407,
   input         cfg_dout1408,
   input         cfg_dout1409,
   input         cfg_dout1410,
   input         cfg_dout1411,
   input         cfg_dout1412,
   input         cfg_dout1413,
   input         cfg_dout1414,
   input         cfg_dout1415,
   input         cfg_dout1416,
   input         cfg_dout1417,
   input         cfg_dout1418,
   input         cfg_dout1419,
   input         cfg_dout1420,
   input         cfg_dout1421,
   input         cfg_dout1422,
   input         cfg_dout1423,
   input         cfg_dout1424,
   input         cfg_dout1425,
   input         cfg_dout1426,
   input         cfg_dout1427,
   input         cfg_dout1428,
   input         cfg_dout1429,
   input         cfg_dout1430,
   input         cfg_dout1431,
   input         cfg_dout1432,
   input         cfg_dout1433,
   input         cfg_dout1434,
   input         cfg_dout1435,
   input         cfg_dout1436,
   input         cfg_dout1437,
   input         cfg_dout1438,
   input         cfg_dout1439,
   input         cfg_dout1440,
   input         cfg_dout1441,
   input         cfg_dout1442,
   input         cfg_dout1443,
   input         cfg_dout1444,
   input         cfg_dout1445,
   input         cfg_dout1446,
   input         cfg_dout1447,
   input         cfg_dout1448,
   input         cfg_dout1449,
   input         cfg_dout1450,
   input         cfg_dout1451,
   input         cfg_dout1452,
   input         cfg_dout1453,
   input         cfg_dout1454,
   input         cfg_dout1455,
   input         cfg_dout1456,
   input         cfg_dout1457,
   input         cfg_dout1458,
   input         cfg_dout1459,
   input         cfg_dout1460,
   input         cfg_dout1461,
   input         cfg_dout1462,
   input         cfg_dout1463,
   input         cfg_dout1464,
   input         cfg_dout1465,
   input         cfg_dout1466,
   input         cfg_dout1467,
   input         cfg_dout1468,
   input         cfg_dout1469,
   input         cfg_dout1470,
   input         cfg_dout1471,
   input         cfg_dout1472,
   input         cfg_dout1473,
   input         cfg_dout1474,
   input         cfg_dout1475,
   input         cfg_dout1476,
   input         cfg_dout1477,
   input         cfg_dout1478,
   input         cfg_dout1479,
   input         cfg_dout1480,
   input         cfg_dout1481,
   input         cfg_dout1482,
   input         cfg_dout1483,
   input         cfg_dout1484,
   input         cfg_dout1485,
   input         cfg_dout1486,
   input         cfg_dout1487,
   input         cfg_dout1488,
   input         cfg_dout1489,
   input         cfg_dout1490,
   input         cfg_dout1491,
   input         cfg_dout1492,
   input         cfg_dout1493,
   input         cfg_dout1494,
   input         cfg_dout1495,
   input         cfg_dout1496,
   input         cfg_dout1497,
   input         cfg_dout1498,
   input         cfg_dout1499,
   input         cfg_dout1500,
   input         cfg_dout1501,
   input         cfg_dout1502,
   input         cfg_dout1503,
   input         cfg_dout1504,
   input         cfg_dout1505,
   input         cfg_dout1506,
   input         cfg_dout1507,
   input         cfg_dout1508,
   input         cfg_dout1509,
   input         cfg_dout1510,
   input         cfg_dout1511,
   input         cfg_dout1512,
   input         cfg_dout1513,
   input         cfg_dout1514,
   input         cfg_dout1515,
   input         cfg_dout1516,
   input         cfg_dout1517,
   input         cfg_dout1518,
   input         cfg_dout1519,
   input         cfg_dout1520,
   input         cfg_dout1521,
   input         cfg_dout1522,
   input         cfg_dout1523,
   input         cfg_dout1524,
   input         cfg_dout1525,
   input         cfg_dout1526,
   input         cfg_dout1527,
   input         cfg_dout1528,
   input         cfg_dout1529,
   input         cfg_dout1530,
   input         cfg_dout1531,
   input         cfg_dout1532,
   input         cfg_dout1533,
   input         cfg_dout1534,
   input         cfg_dout1535,
   input         cfg_dout1536,
   input         cfg_dout1537,
   input         cfg_dout1538,
   input         cfg_dout1539,
   input         cfg_dout1540,
   input         cfg_dout1541,
   input         cfg_dout1542,
   input         cfg_dout1543,
   input         cfg_dout1544,
   input         cfg_dout1545,
   input         cfg_dout1546,
   input         cfg_dout1547,
   input         cfg_dout1548,
   input         cfg_dout1549,
   input         cfg_dout1550,
   input         cfg_dout1551,
   input         cfg_dout1552,
   input         cfg_dout1553,
   input         cfg_dout1554,
   input         cfg_dout1555,
   input         cfg_dout1556,
   input         cfg_dout1557,
   input         cfg_dout1558,
   input         cfg_dout1559,
   input         cfg_dout1560,
   input         cfg_dout1561,
   input         cfg_dout1562,
   input         cfg_dout1563,
   input         cfg_dout1564,
   input         cfg_dout1565,
   input         cfg_dout1566,
   input         cfg_dout1567,
   input         cfg_dout1568,
   input         cfg_dout1569,
   input         cfg_dout1570,
   input         cfg_dout1571,
   input         cfg_dout1572,
   input         cfg_dout1573,
   input         cfg_dout1574,
   input         cfg_dout1575,
   input         cfg_dout1576,
   input         cfg_dout1577,
   input         cfg_dout1578,
   input         cfg_dout1579,
   input         cfg_dout1580,
   input         cfg_dout1581,
   input         cfg_dout1582,
   input         cfg_dout1583,
   input         cfg_dout1584,
   input         cfg_dout1585,
   input         cfg_dout1586,
   input         cfg_dout1587,
   input         cfg_dout1588,
   input         cfg_dout1589,
   input         cfg_dout1590,
   input         cfg_dout1591,
   input         cfg_dout1592,
   input         cfg_dout1593,
   input         cfg_dout1594,
   input         cfg_dout1595,
   input         cfg_dout1596,
   input         cfg_dout1597,
   input         cfg_dout1598,
   input         cfg_dout1599,
   input         cfg_dout1600,
   input         cfg_dout1601,
   input         cfg_dout1602,
   input         cfg_dout1603,
   input         cfg_dout1604,
   input         cfg_dout1605,
   input         cfg_dout1606,
   input         cfg_dout1607,
   input         cfg_dout1608,
   input         cfg_dout1609,
   input         cfg_dout1610,
   input         cfg_dout1611,
   input         cfg_dout1612,
   input         cfg_dout1613,
   input         cfg_dout1614,
   input         cfg_dout1615,
   input         cfg_dout1616,
   input         cfg_dout1617,
   input         cfg_dout1618,
   input         cfg_dout1619,
   input         cfg_dout1620,
   input         cfg_dout1621,
   input         cfg_dout1622,
   input         cfg_dout1623,
   input         cfg_dout1624,
   input         cfg_dout1625,
   input         cfg_dout1626,
   input         cfg_dout1627,
   input         cfg_dout1628,
   input         cfg_dout1629,
   input         cfg_dout1630,
   input         cfg_dout1631,
   input         cfg_dout1632,
   input         cfg_dout1633,
   input         cfg_dout1634,
   input         cfg_dout1635,
   input         cfg_dout1636,
   input         cfg_dout1637,
   input         cfg_dout1638,
   input         cfg_dout1639,
   input         cfg_dout1640,
   input         cfg_dout1641,
   input         cfg_dout1642,
   input         cfg_dout1643,
   input         cfg_dout1644,
   input         cfg_dout1645,
   input         cfg_dout1646,
   input         cfg_dout1647,
   input         cfg_dout1648,
   input         cfg_dout1649,
   input         cfg_dout1650,
   input         cfg_dout1651,
   input         cfg_dout1652,
   input         cfg_dout1653,
   input         cfg_dout1654,
   input         cfg_dout1655,
   input         cfg_dout1656,
   input         cfg_dout1657,
   input         cfg_dout1658,
   input         cfg_dout1659,
   input         cfg_dout1660,
   input         cfg_dout1661,
   input         cfg_dout1662,
   input         cfg_dout1663,
   input         cfg_dout1664,
   input         cfg_dout1665,
   input         cfg_dout1666,
   input         cfg_dout1667,
   input         cfg_dout1668,
   input         cfg_dout1669,
   input         cfg_dout1670,
   input         cfg_dout1671,
   input         cfg_dout1672,
   input         cfg_dout1673,
   input         cfg_dout1674,
   input         cfg_dout1675,
   input         cfg_dout1676,
   input         cfg_dout1677,
   input         cfg_dout1678,
   input         cfg_dout1679,
   input         cfg_dout1680,
   input         cfg_dout1681,
   input         cfg_dout1682,
   input         cfg_dout1683,
   input         cfg_dout1684,
   input         cfg_dout1685,
   input         cfg_dout1686,
   input         cfg_dout1687,
   input         cfg_dout1688,
   input         cfg_dout1689,
   input         cfg_dout1690,
   input         cfg_dout1691,
   input         cfg_dout1692,
   input         cfg_dout1693,
   input         cfg_dout1694,
   input         cfg_dout1695,
   input         cfg_dout1696,
   input         cfg_dout1697,
   input         cfg_dout1698,
   input         cfg_dout1699,
   input         cfg_dout1700,
   input         cfg_dout1701,
   input         cfg_dout1702,
   input         cfg_dout1703,
   input         cfg_dout1704,
   input         cfg_dout1705,
   input         cfg_dout1706,
   input         cfg_dout1707,
   input         cfg_dout1708,
   input         cfg_dout1709,
   input         cfg_dout1710,
   input         cfg_dout1711,
   input         cfg_dout1712,
   input         cfg_dout1713,
   input         cfg_dout1714,
   input         cfg_dout1715,
   input         cfg_dout1716,
   input         cfg_dout1717,
   input         cfg_dout1718,
   input         cfg_dout1719,
   input         cfg_dout1720,
   input         cfg_dout1721,
   input         cfg_dout1722,
   input         cfg_dout1723,
   input         cfg_dout1724,
   input         cfg_dout1725,
   input         cfg_dout1726,
   input         cfg_dout1727,
   input         cfg_dout1728,
   input         cfg_dout1729,
   input         cfg_dout1730,
   input         cfg_dout1731,
   input         cfg_dout1732,
   input         cfg_dout1733,
   input         cfg_dout1734,
   input         cfg_dout1735,
   input         cfg_dout1736,
   input         cfg_dout1737,
   input         cfg_dout1738,
   input         cfg_dout1739,
   input         cfg_dout1740,
   input         cfg_dout1741,
   input         cfg_dout1742,
   input         cfg_dout1743,
   input         cfg_dout1744,
   input         cfg_dout1745,
   input         cfg_dout1746,
   input         cfg_dout1747,
   input         cfg_dout1748,
   input         cfg_dout1749,
   input         cfg_dout1750,
   input         cfg_dout1751,
   input         cfg_dout1752,
   input         cfg_dout1753,
   input         cfg_dout1754,
   input         cfg_dout1755,
   input         cfg_dout1756,
   input         cfg_dout1757,
   input         cfg_dout1758,
   input         cfg_dout1759,
   input         cfg_dout1760,
   input         cfg_dout1761,
   input         cfg_dout1762,
   input         cfg_dout1763,
   input         cfg_dout1764,
   input         cfg_dout1765,
   input         cfg_dout1766,
   input         cfg_dout1767,
   input         cfg_dout1768,
   input         cfg_dout1769,
   input         cfg_dout1770,
   input         cfg_dout1771,
   input         cfg_dout1772,
   input         cfg_dout1773,
   input         cfg_dout1774,
   input         cfg_dout1775,
   input         cfg_dout1776,
   input         cfg_dout1777,
   input         cfg_dout1778,
   input         cfg_dout1779,
   input         cfg_dout1780,
   input         cfg_dout1781,
   input         cfg_dout1782,
   input         cfg_dout1783,
   input         cfg_dout1784,
   input         cfg_dout1785,
   input         cfg_dout1786,
   input         cfg_dout1787,
   input         cfg_dout1788,
   input         cfg_dout1789,
   input         cfg_dout1790,
   input         cfg_dout1791,
   input         cfg_dout1792,
   input         cfg_dout1793,
   input         cfg_dout1794,
   input         cfg_dout1795,
   input         cfg_dout1796,
   input         cfg_dout1797,
   input         cfg_dout1798,
   input         cfg_dout1799,
   input         cfg_dout1800,
   input         cfg_dout1801,
   input         cfg_dout1802,
   input         cfg_dout1803,
   input         cfg_dout1804,
   input         cfg_dout1805,
   input         cfg_dout1806,
   input         cfg_dout1807,
   input         cfg_dout1808,
   input         cfg_dout1809,
   input         cfg_dout1810,
   input         cfg_dout1811,
   input         cfg_dout1812,
   input         cfg_dout1813,
   input         cfg_dout1814,
   input         cfg_dout1815,
   input         cfg_dout1816,
   input         cfg_dout1817,
   input         cfg_dout1818,
   input         cfg_dout1819,
   input         cfg_dout1820,
   input         cfg_dout1821,
   input         cfg_dout1822,
   input         cfg_dout1823,
   input         cfg_dout1824,
   input         cfg_dout1825,
   input         cfg_dout1826,
   input         cfg_dout1827,
   input         cfg_dout1828,
   input         cfg_dout1829,
   input         cfg_dout1830,
   input         cfg_dout1831,
   input         cfg_dout1832,
   input         cfg_dout1833,
   input         cfg_dout1834,
   input         cfg_dout1835,
   input         cfg_dout1836,
   input         cfg_dout1837,
   input         cfg_dout1838,
   input         cfg_dout1839,
   input         cfg_dout1840,
   input         cfg_dout1841,
   input         cfg_dout1842,
   input         cfg_dout1843,
   input         cfg_dout1844,
   input         cfg_dout1845,
   input         cfg_dout1846,
   input         cfg_dout1847,
   input         cfg_dout1848,
   input         cfg_dout1849,
   input         cfg_dout1850,
   input         cfg_dout1851,
   input         cfg_dout1852,
   input         cfg_dout1853,
   input         cfg_dout1854,
   input         cfg_dout1855,
   input         cfg_dout1856,
   input         cfg_dout1857,
   input         cfg_dout1858,
   input         cfg_dout1859,
   input         cfg_dout1860,
   input         cfg_dout1861,
   input         cfg_dout1862,
   input         cfg_dout1863,
   input         cfg_dout1864,
   input         cfg_dout1865,
   input         cfg_dout1866,
   input         cfg_dout1867,
   input         cfg_dout1868,
   input         cfg_dout1869,
   input         cfg_dout1870,
   input         cfg_dout1871,
   input         cfg_dout1872,
   input         cfg_dout1873,
   input         cfg_dout1874,
   input         cfg_dout1875,
   input         cfg_dout1876,
   input         cfg_dout1877,
   input         cfg_dout1878,
   input         cfg_dout1879,
   input         cfg_dout1880,
   input         cfg_dout1881,
   input         cfg_dout1882,
   input         cfg_dout1883,
   input         cfg_dout1884,
   input         cfg_dout1885,
   input         cfg_dout1886,
   input         cfg_dout1887,
   input         cfg_dout1888,
   input         cfg_dout1889,
   input         cfg_dout1890,
   input         cfg_dout1891,
   input         cfg_dout1892,
   input         cfg_dout1893,
   input         cfg_dout1894,
   input         cfg_dout1895,
   input         cfg_dout1896,
   input         cfg_dout1897,
   input         cfg_dout1898,
   input         cfg_dout1899,
   input         cfg_dout1900,
   input         cfg_dout1901,
   input         cfg_dout1902,
   input         cfg_dout1903,
   input         cfg_dout1904,
   input         cfg_dout1905,
   input         cfg_dout1906,
   input         cfg_dout1907,
   input         cfg_dout1908,
   input         cfg_dout1909,
   input         cfg_dout1910,
   input         cfg_dout1911,
   input         cfg_dout1912,
   input         cfg_dout1913,
   input         cfg_dout1914,
   input         cfg_dout1915,
   input         cfg_dout1916,
   input         cfg_dout1917,
   input         cfg_dout1918,
   input         cfg_dout1919,
   input         cfg_dout1920,
   input         cfg_dout1921,
   input         cfg_dout1922,
   input         cfg_dout1923,
   input         cfg_dout1924,
   input         cfg_dout1925,
   input         cfg_dout1926,
   input         cfg_dout1927,
   input         cfg_dout1928,
   input         cfg_dout1929,
   input         cfg_dout1930,
   input         cfg_dout1931,
   input         cfg_dout1932,
   input         cfg_dout1933,
   input         cfg_dout1934,
   input         cfg_dout1935,
   input         cfg_dout1936,
   input         cfg_dout1937,
   input         cfg_dout1938,
   input         cfg_dout1939,
   input         cfg_dout1940,
   input         cfg_dout1941,
   input         cfg_dout1942,
   input         cfg_dout1943,
   input         cfg_dout1944,
   input         cfg_dout1945,
   input         cfg_dout1946,
   input         cfg_dout1947,
   input         cfg_dout1948,
   input         cfg_dout1949,
   input         cfg_dout1950,
   input         cfg_dout1951,
   input         cfg_dout1952,
   input         cfg_dout1953,
   input         cfg_dout1954,
   input         cfg_dout1955,
   input         cfg_dout1956,
   input         cfg_dout1957,
   input         cfg_dout1958,
   input         cfg_dout1959,
   input         cfg_dout1960,
   input         cfg_dout1961,
   input         cfg_dout1962,
   input         cfg_dout1963,
   input         cfg_dout1964,
   input         cfg_dout1965,
   input         cfg_dout1966,
   input         cfg_dout1967,
   input         cfg_dout1968,
   input         cfg_dout1969,
   input         cfg_dout1970,
   input         cfg_dout1971,
   input         cfg_dout1972,
   input         cfg_dout1973,
   input         cfg_dout1974,
   input         cfg_dout1975,
   input         cfg_dout1976,
   input         cfg_dout1977,
   input         cfg_dout1978,
   input         cfg_dout1979,
   input         cfg_dout1980,
   input         cfg_dout1981,
   input         cfg_dout1982,
   input         cfg_dout1983,
   input         cfg_dout1984,
   input         cfg_dout1985,
   input         cfg_dout1986,
   input         cfg_dout1987,
   input         cfg_dout1988,
   input         cfg_dout1989,
   input         cfg_dout1990,
   input         cfg_dout1991,
   input         cfg_dout1992,
   input         cfg_dout1993,
   input         cfg_dout1994,
   input         cfg_dout1995,
   input         cfg_dout1996,
   input         cfg_dout1997,
   input         cfg_dout1998,
   input         cfg_dout1999,
   input         cfg_dout2000,
   input         cfg_dout2001,
   input         cfg_dout2002,
   input         cfg_dout2003,
   input         cfg_dout2004,
   input         cfg_dout2005,
   input         cfg_dout2006,
   input         cfg_dout2007,
   input         cfg_dout2008,
   input         cfg_dout2009,
   input         cfg_dout2010,
   input         cfg_dout2011,
   input         cfg_dout2012,
   input         cfg_dout2013,
   input         cfg_dout2014,
   input         cfg_dout2015,
   input         cfg_dout2016,
   input         cfg_dout2017,
   input         cfg_dout2018,
   input         cfg_dout2019,
   input         cfg_dout2020,
   input         cfg_dout2021,
   input         cfg_dout2022,
   input         cfg_dout2023,
   input         cfg_dout2024,
   input         cfg_dout2025,
   input         cfg_dout2026,
   input         cfg_dout2027,
   input         cfg_dout2028,
   input         cfg_dout2029,
   input         cfg_dout2030,
   input         cfg_dout2031,
   input         cfg_dout2032,
   input         cfg_dout2033,
   input         cfg_dout2034,
   input         cfg_dout2035,
   input         cfg_dout2036,
   input         cfg_dout2037,
   input         cfg_dout2038,
   input         cfg_dout2039,
   input         cfg_dout2040,
   input         cfg_dout2041,
   input         cfg_dout2042,
   input         cfg_dout2043,
   input         cfg_dout2044,
   input         cfg_dout2045,
   input         cfg_dout2046,
   input         cfg_dout2047,
   input         cfg_dout2048,
   input         cfg_dout2049,
   input         cfg_dout2050,
   input         cfg_dout2051,
   input         cfg_dout2052,
   input         cfg_dout2053,
   input         cfg_dout2054,
   input         cfg_dout2055,
   input         cfg_dout2056,
   input         cfg_dout2057,
   input         cfg_dout2058,
   input         cfg_dout2059,
   input         cfg_dout2060,
   input         cfg_dout2061,
   input         cfg_dout2062,
   input         cfg_dout2063,
   input         cfg_dout2064,
   input         cfg_dout2065,
   input         cfg_dout2066,
   input         cfg_dout2067,
   input         cfg_dout2068,
   input         cfg_dout2069,
   input         cfg_dout2070,
   input         cfg_dout2071,
   input         cfg_dout2072,
   input         cfg_dout2073,
   input         cfg_dout2074,
   input         cfg_dout2075,
   input         cfg_dout2076,
   input         cfg_dout2077,
   input         cfg_dout2078,
   input         cfg_dout2079,
   input         cfg_dout2080,
   input         cfg_dout2081,
   input         cfg_dout2082,
   input         cfg_dout2083,
   input         cfg_dout2084,
   input         cfg_dout2085,
   input         cfg_dout2086,
   input         cfg_dout2087,
   input         cfg_dout2088,
   input         cfg_dout2089,
   input         cfg_dout2090,
   input         cfg_dout2091,
   input         cfg_dout2092,
   input         cfg_dout2093,
   input         cfg_dout2094,
   input         cfg_dout2095,
   input         cfg_dout2096,
   input         cfg_dout2097,
   input         cfg_dout2098,
   input         cfg_dout2099,
   input         cfg_dout2100,
   input         cfg_dout2101,
   input         cfg_dout2102,
   input         cfg_dout2103,
   input         cfg_dout2104,
   input         cfg_dout2105,
   input         cfg_dout2106,
   input         cfg_dout2107,
   input         cfg_dout2108,
   input         cfg_dout2109,
   input         cfg_dout2110,
   input         cfg_dout2111,
   input         cfg_dout2112,
   input         cfg_dout2113,
   input         cfg_dout2114,
   input         cfg_dout2115,
   input         cfg_dout2116,
   input         cfg_dout2117,
   input         cfg_dout2118,
   input         cfg_dout2119,
   input         cfg_dout2120,
   input         cfg_dout2121,
   input         cfg_dout2122,
   input         cfg_dout2123,
   input         cfg_dout2124,
   input         cfg_dout2125,
   input         cfg_dout2126,
   input         cfg_dout2127,
   input         cfg_dout2128,
   input         cfg_dout2129,
   input         cfg_dout2130,
   input         cfg_dout2131,
   input         cfg_dout2132,
   input         cfg_dout2133,
   input         cfg_dout2134,
   input         cfg_dout2135,
   input         cfg_dout2136,
   input         cfg_dout2137,
   input         cfg_dout2138,
   input         cfg_dout2139,
   input         cfg_dout2140,
   input         cfg_dout2141,
   input         cfg_dout2142,
   input         cfg_dout2143,
   input         cfg_dout2144,
   input         cfg_dout2145,
   input         cfg_dout2146,
   input         cfg_dout2147,
   input         cfg_dout2148,
   input         cfg_dout2149,
   input         cfg_dout2150,
   input         cfg_dout2151,
   input         cfg_dout2152,
   input         cfg_dout2153,
   input         cfg_dout2154,
   input         cfg_dout2155,
   input         cfg_dout2156,
   input         cfg_dout2157,
   input         cfg_dout2158,
   input         cfg_dout2159,
   input         cfg_dout2160,
   input         cfg_dout2161,
   input         cfg_dout2162,
   input         cfg_dout2163,
   input         cfg_dout2164,
   input         cfg_dout2165,
   input         cfg_dout2166,
   input         cfg_dout2167,
   input         cfg_dout2168,
   input         cfg_dout2169,
   input         cfg_dout2170,
   input         cfg_dout2171,
   input         cfg_dout2172,
   input         cfg_dout2173,
   input         cfg_dout2174,
   input         cfg_dout2175,
   input         cfg_dout2176,
   input         cfg_dout2177,
   input         cfg_dout2178,
   input         cfg_dout2179,
   input         cfg_dout2180,
   input         cfg_dout2181,
   input         cfg_dout2182,
   input         cfg_dout2183,
   input         cfg_dout2184,
   input         cfg_dout2185,
   input         cfg_dout2186,
   input         cfg_dout2187,
   input         cfg_dout2188,
   input         cfg_dout2189,
   input         cfg_dout2190,
   input         cfg_dout2191,
   input         cfg_dout2192,
   input         cfg_dout2193,
   input         cfg_dout2194,
   input         cfg_dout2195,
   input         cfg_dout2196,
   input         cfg_dout2197,
   input         cfg_dout2198,
   input         cfg_dout2199,
   input         cfg_dout2200,
   input         cfg_dout2201,
   input         cfg_dout2202,
   input         cfg_dout2203,
   input         cfg_dout2204,
   input         cfg_dout2205,
   input         cfg_dout2206,
   input         cfg_dout2207,
   input         cfg_dout2208,
   input         cfg_dout2209,
   input         cfg_dout2210,
   input         cfg_dout2211,
   input         cfg_dout2212,
   input         cfg_dout2213,
   input         cfg_dout2214,
   input         cfg_dout2215,
   input         cfg_dout2216,
   input         cfg_dout2217,
   input         cfg_dout2218,
   input         cfg_dout2219,
   input         cfg_dout2220,
   input         cfg_dout2221,
   input         cfg_dout2222,
   input         cfg_dout2223,
   input         cfg_dout2224,
   input         cfg_dout2225,
   input         cfg_dout2226,
   input         cfg_dout2227,
   input         cfg_dout2228,
   input         cfg_dout2229,
   input         cfg_dout2230,
   input         cfg_dout2231,
   input         cfg_dout2232,
   input         cfg_dout2233,
   input         cfg_dout2234,
   input         cfg_dout2235,
   input         cfg_dout2236,
   input         cfg_dout2237,
   input         cfg_dout2238,
   input         cfg_dout2239,
   input         cfg_dout2240,
   input         cfg_dout2241,
   input         cfg_dout2242,
   input         cfg_dout2243,
   input         cfg_dout2244,
   input         cfg_dout2245,
   input         cfg_dout2246,
   input         cfg_dout2247,
   input         cfg_dout2248,
   input         cfg_dout2249,
   input         cfg_dout2250,
   input         cfg_dout2251,
   input         cfg_dout2252,
   input         cfg_dout2253,
   input         cfg_dout2254,
   input         cfg_dout2255,
   input         cfg_dout2256,
   input         cfg_dout2257,
   input         cfg_dout2258,
   input         cfg_dout2259,
   input         cfg_dout2260,
   input         cfg_dout2261,
   input         cfg_dout2262,
   input         cfg_dout2263,
   input         cfg_dout2264,
   input         cfg_dout2265,
   input         cfg_dout2266,
   input         cfg_dout2267,
   input         cfg_dout2268,
   input         cfg_dout2269,
   input         cfg_dout2270,
   input         cfg_dout2271,
   input         cfg_dout2272,
   input         cfg_dout2273,
   input         cfg_dout2274,
   input         cfg_dout2275,
   input         cfg_dout2276,
   input         cfg_dout2277,
   input         cfg_dout2278,
   input         cfg_dout2279,
   input         cfg_dout2280,
   input         cfg_dout2281,
   input         cfg_dout2282,
   input         cfg_dout2283,
   input         cfg_dout2284,
   input         cfg_dout2285,
   input         cfg_dout2286,
   input         cfg_dout2287,
   input         cfg_dout2288,
   input         cfg_dout2289,
   input         cfg_dout2290,
   input         cfg_dout2291,
   input         cfg_dout2292,
   input         cfg_dout2293,
   input         cfg_dout2294,
   input         cfg_dout2295,
   input         cfg_dout2296,
   input         cfg_dout2297,
   input         cfg_dout2298,
   input         cfg_dout2299,
   input         cfg_dout2300,
   input         cfg_dout2301,
   input         cfg_dout2302,
   input         cfg_dout2303,
   input         cfg_dout2304,
   input         cfg_dout2305,
   input         cfg_dout2306,
   input         cfg_dout2307,
   input         cfg_dout2308,
   input         cfg_dout2309,
   input         cfg_dout2310,
   input         cfg_dout2311,
   input         cfg_dout2312,
   input         cfg_dout2313,
   input         cfg_dout2314,
   input         cfg_dout2315,
   input         cfg_dout2316,
   input         cfg_dout2317,
   input         cfg_dout2318,
   input         cfg_dout2319,
   input         cfg_dout2320,
   input         cfg_dout2321,
   input         cfg_dout2322,
   input         cfg_dout2323,
   input         cfg_dout2324,
   input         cfg_dout2325,
   input         cfg_dout2326,
   input         cfg_dout2327,
   input         cfg_dout2328,
   input         cfg_dout2329,
   input         cfg_dout2330,
   input         cfg_dout2331,
   input         cfg_dout2332,
   input         cfg_dout2333,
   input         cfg_dout2334,
   input         cfg_dout2335,
   input         cfg_dout2336,
   input         cfg_dout2337,
   input         cfg_dout2338,
   input         cfg_dout2339,
   input         cfg_dout2340,
   input         cfg_dout2341,
   input         cfg_dout2342,
   input         cfg_dout2343,
   input         cfg_dout2344,
   input         cfg_dout2345,
   input         cfg_dout2346,
   input         cfg_dout2347,
   input         cfg_dout2348,
   input         cfg_dout2349,
   input         cfg_dout2350,
   input         cfg_dout2351,
   input         cfg_dout2352,
   input         cfg_dout2353,
   input         cfg_dout2354,
   input         cfg_dout2355,
   input         cfg_dout2356,
   input         cfg_dout2357,
   input         cfg_dout2358,
   input         cfg_dout2359,
   input         cfg_dout2360,
   input         cfg_dout2361,
   input         cfg_dout2362,
   input         cfg_dout2363,
   input         cfg_dout2364,
   input         cfg_dout2365,
   input         cfg_dout2366,
   input         cfg_dout2367,
   input         cfg_dout2368,
   input         cfg_dout2369,
   input         cfg_dout2370,
   input         cfg_dout2371,
   input         cfg_dout2372,
   input         cfg_dout2373,
   input         cfg_dout2374,
   input         cfg_dout2375,
   input         cfg_dout2376,
   input         cfg_dout2377,
   input         cfg_dout2378,
   input         cfg_dout2379,
   input         cfg_dout2380,
   input         cfg_dout2381,
   input         cfg_dout2382,
   input         cfg_dout2383,
   input         cfg_dout2384,
   input         cfg_dout2385,
   input         cfg_dout2386,
   input         cfg_dout2387,
   input         cfg_dout2388,
   input         cfg_dout2389,
   input         cfg_dout2390,
   input         cfg_dout2391,
   input         cfg_dout2392,
   input         cfg_dout2393,
   input         cfg_dout2394,
   input         cfg_dout2395,
   input         cfg_dout2396,
   input         cfg_dout2397,
   input         cfg_dout2398,
   input         cfg_dout2399,
   input         cfg_dout2400,
   input         cfg_dout2401,
   input         cfg_dout2402,
   input         cfg_dout2403,
   input         cfg_dout2404,
   input         cfg_dout2405,
   input         cfg_dout2406,
   input         cfg_dout2407,
   input         cfg_dout2408,
   input         cfg_dout2409,
   input         cfg_dout2410,
   input         cfg_dout2411,
   input         cfg_dout2412,
   input         cfg_dout2413,
   input         cfg_dout2414,
   input         cfg_dout2415,
   input         cfg_dout2416,
   input         cfg_dout2417,
   input         cfg_dout2418,
   input         cfg_dout2419,
   input         cfg_dout2420,
   input         cfg_dout2421,
   input         cfg_dout2422,
   input         cfg_dout2423,
   input         cfg_dout2424,
   input         cfg_dout2425,
   input         cfg_dout2426,
   input         cfg_dout2427,
   input         cfg_dout2428,
   input         cfg_dout2429,
   input         cfg_dout2430,
   input         cfg_dout2431,
   input         cfg_dout2432,
   input         cfg_dout2433,
   input         cfg_dout2434,
   input         cfg_dout2435,
   input         cfg_dout2436,
   input         cfg_dout2437,
   input         cfg_dout2438,
   input         cfg_dout2439,
   input         cfg_dout2440,
   input         cfg_dout2441,
   input         cfg_dout2442,
   input         cfg_dout2443,
   input         cfg_dout2444,
   input         cfg_dout2445,
   input         cfg_dout2446,
   input         cfg_dout2447,
   input         cfg_dout2448,
   input         cfg_dout2449,
   input         cfg_dout2450,
   input         cfg_dout2451,
   input         cfg_dout2452,
   input         cfg_dout2453,
   input         cfg_dout2454,
   input         cfg_dout2455,
   input         cfg_dout2456,
   input         cfg_dout2457,
   input         cfg_dout2458,
   input         cfg_dout2459,
   input         cfg_dout2460,
   input         cfg_dout2461,
   input         cfg_dout2462,
   input         cfg_dout2463,
   input         cfg_dout2464,
   input         cfg_dout2465,
   input         cfg_dout2466,
   input         cfg_dout2467,
   input         cfg_dout2468,
   input         cfg_dout2469,
   input         cfg_dout2470,
   input         cfg_dout2471,
   input         cfg_dout2472,
   input         cfg_dout2473,
   input         cfg_dout2474,
   input         cfg_dout2475,
   input         cfg_dout2476,
   input         cfg_dout2477,
   input         cfg_dout2478,
   input         cfg_dout2479,
   input         cfg_dout2480,
   input         cfg_dout2481,
   input         cfg_dout2482,
   input         cfg_dout2483,
   input         cfg_dout2484,
   input         cfg_dout2485,
   input         cfg_dout2486,
   input         cfg_dout2487,
   input         cfg_dout2488,
   input         cfg_dout2489,
   input         cfg_dout2490,
   input         cfg_dout2491,
   input         cfg_dout2492,
   input         cfg_dout2493,
   input         cfg_dout2494,
   input         cfg_dout2495,
   input         cfg_dout2496,
   input         cfg_dout2497,
   input         cfg_dout2498,
   input         cfg_dout2499,
   input         cfg_dout2500,
   input         cfg_dout2501,
   input         cfg_dout2502,
   input         cfg_dout2503,
   input         cfg_dout2504,
   input         cfg_dout2505,
   input         cfg_dout2506,
   input         cfg_dout2507,
   input         cfg_dout2508,
   input         cfg_dout2509,
   input         cfg_dout2510,
   input         cfg_dout2511,
   input         cfg_dout2512,
   input         cfg_dout2513,
   input         cfg_dout2514,
   input         cfg_dout2515,
   input         cfg_dout2516,
   input         cfg_dout2517,
   input         cfg_dout2518,
   input         cfg_dout2519,
   input         cfg_dout2520,
   input         cfg_dout2521,
   input         cfg_dout2522,
   input         cfg_dout2523,
   input         cfg_dout2524,
   input         cfg_dout2525,
   input         cfg_dout2526,
   input         cfg_dout2527,
   input         cfg_dout2528,
   input         cfg_dout2529,
   input         cfg_dout2530,
   input         cfg_dout2531,
   input         cfg_dout2532,
   input         cfg_dout2533,
   input         cfg_dout2534,
   input         cfg_dout2535,
   input         cfg_dout2536,
   input         cfg_dout2537,
   input         cfg_dout2538,
   input         cfg_dout2539,
   input         cfg_dout2540,
   input         cfg_dout2541,
   input         cfg_dout2542,
   input         cfg_dout2543,
   input         cfg_dout2544,
   input         cfg_dout2545,
   input         cfg_dout2546,
   input         cfg_dout2547,
   input         cfg_dout2548,
   input         cfg_dout2549,
   input         cfg_dout2550,
   input         cfg_dout2551,
   input         cfg_dout2552,
   input         cfg_dout2553,
   input         cfg_dout2554,
   input         cfg_dout2555,
   input         cfg_dout2556,
   input         cfg_dout2557,
   input         cfg_dout2558,
   input         cfg_dout2559,
   input         cfg_dout2560,
   input         cfg_dout2561,
   input         cfg_dout2562,
   input         cfg_dout2563,
   input         cfg_dout2564,
   input         cfg_dout2565,
   input         cfg_dout2566,
   input         cfg_dout2567,
   input         cfg_dout2568,
   input         cfg_dout2569,
   input         cfg_dout2570,
   input         cfg_dout2571,
   input         cfg_dout2572,
   input         cfg_dout2573,
   input         cfg_dout2574,
   input         cfg_dout2575,
   input         cfg_dout2576,
   input         cfg_dout2577,
   input         cfg_dout2578,
   input         cfg_dout2579,
   input         cfg_dout2580,
   input         cfg_dout2581,
   input         cfg_dout2582,
   input         cfg_dout2583,
   input         cfg_dout2584,
   input         cfg_dout2585,
   input         cfg_dout2586,
   input         cfg_dout2587,
   input         cfg_dout2588,
   input         cfg_dout2589,
   input         cfg_dout2590,
   input         cfg_dout2591,
   input         cfg_dout2592,
   input         cfg_dout2593,
   input         cfg_dout2594,
   input         cfg_dout2595,
   input         cfg_dout2596,
   input         cfg_dout2597,
   input         cfg_dout2598,
   input         cfg_dout2599,
   input         cfg_dout2600,
   input         cfg_dout2601,
   input         cfg_dout2602,
   input         cfg_dout2603,
   input         cfg_dout2604,
   input         cfg_dout2605,
   input         cfg_dout2606,
   input         cfg_dout2607,
   input         cfg_dout2608,
   input         cfg_dout2609,
   input         cfg_dout2610,
   input         cfg_dout2611,
   input         cfg_dout2612,
   input         cfg_dout2613,
   input         cfg_dout2614,
   input         cfg_dout2615,
   input         cfg_dout2616,
   input         cfg_dout2617,
   input         cfg_dout2618,
   input         cfg_dout2619,
   input         cfg_dout2620,
   input         cfg_dout2621,
   input         cfg_dout2622,
   input         cfg_dout2623,
   input         cfg_dout2624,
   input         cfg_dout2625,
   input         cfg_dout2626,
   input         cfg_dout2627,
   input         cfg_dout2628,
   input         cfg_dout2629,
   input         cfg_dout2630,
   input         cfg_dout2631,
   input         cfg_dout2632,
   input         cfg_dout2633,
   input         cfg_dout2634,
   input         cfg_dout2635,
   input         cfg_dout2636,
   input         cfg_dout2637,
   input         cfg_dout2638,
   input         cfg_dout2639,
   input         cfg_dout2640,
   input         cfg_dout2641,
   input         cfg_dout2642,
   input         cfg_dout2643,
   input         cfg_dout2644,
   input         cfg_dout2645,
   input         cfg_dout2646,
   input         cfg_dout2647,
   input         cfg_dout2648,
   input         cfg_dout2649,
   input         cfg_dout2650,
   input         cfg_dout2651,
   input         cfg_dout2652,
   input         cfg_dout2653,
   input         cfg_dout2654,
   input         cfg_dout2655,
   input         cfg_dout2656,
   input         cfg_dout2657,
   input         cfg_dout2658,
   input         cfg_dout2659,
   input         cfg_dout2660,
   input         cfg_dout2661,
   input         cfg_dout2662,
   input         cfg_dout2663,
   input         cfg_dout2664,
   input         cfg_dout2665,
   input         cfg_dout2666,
   input         cfg_dout2667,
   input         cfg_dout2668,
   input         cfg_dout2669,
   input         cfg_dout2670,
   input         cfg_dout2671,
   input         cfg_dout2672,
   input         cfg_dout2673,
   input         cfg_dout2674,
   input         cfg_dout2675,
   input         cfg_dout2676,
   input         cfg_dout2677,
   input         cfg_dout2678,
   input         cfg_dout2679,
   input         cfg_dout2680,
   input         cfg_dout2681,
   input         cfg_dout2682,
   input         cfg_dout2683,
   input         cfg_dout2684,
   input         cfg_dout2685,
   input         cfg_dout2686,
   input         cfg_dout2687,
   input         cfg_dout2688,
   input         cfg_dout2689,
   input         cfg_dout2690,
   input         cfg_dout2691,
   input         cfg_dout2692,
   input         cfg_dout2693,
   input         cfg_dout2694,
   input         cfg_dout2695,
   input         cfg_dout2696,
   input         cfg_dout2697,
   input         cfg_dout2698,
   input         cfg_dout2699,
   input         cfg_dout2700,
   input         cfg_dout2701,
   input         cfg_dout2702,
   input         cfg_dout2703,
   input         cfg_dout2704,
   input         cfg_dout2705,
   input         cfg_dout2706,
   input         cfg_dout2707,
   input         cfg_dout2708,
   input         cfg_dout2709,
   input         cfg_dout2710,
   input         cfg_dout2711,
   input         cfg_dout2712,
   input         cfg_dout2713,
   input         cfg_dout2714,
   input         cfg_dout2715,
   input         cfg_dout2716,
   input         cfg_dout2717,
   input         cfg_dout2718,
   input         cfg_dout2719,
   input         cfg_dout2720,
   input         cfg_dout2721,
   input         cfg_dout2722,
   input         cfg_dout2723,
   input         cfg_dout2724,
   input         cfg_dout2725,
   input         cfg_dout2726,
   input         cfg_dout2727,
   input         cfg_dout2728,
   input         cfg_dout2729,
   input         cfg_dout2730,
   input         cfg_dout2731,
   input         cfg_dout2732,
   input         cfg_dout2733,
   input         cfg_dout2734,
   input         cfg_dout2735,
   input         cfg_dout2736,
   input         cfg_dout2737,
   input         cfg_dout2738,
   input         cfg_dout2739,
   input         cfg_dout2740,
   input         cfg_dout2741,
   input         cfg_dout2742,
   input         cfg_dout2743,
   input         cfg_dout2744,
   input         cfg_dout2745,
   input         cfg_dout2746,
   input         cfg_dout2747,
   input         cfg_dout2748,
   input         cfg_dout2749,
   input         cfg_dout2750,
   input         cfg_dout2751,
   input         cfg_dout2752,
   input         cfg_dout2753,
   input         cfg_dout2754,
   input         cfg_dout2755,
   input         cfg_dout2756,
   input         cfg_dout2757,
   input         cfg_dout2758,
   input         cfg_dout2759,
   input         cfg_dout2760,
   input         cfg_dout2761,
   input         cfg_dout2762,
   input         cfg_dout2763,
   input         cfg_dout2764,
   input         cfg_dout2765,
   input         cfg_dout2766,
   input         cfg_dout2767,
   input         cfg_dout2768,
   input         cfg_dout2769,
   input         cfg_dout2770,
   input         cfg_dout2771,
   input         cfg_dout2772,
   input         cfg_dout2773,
   input         cfg_dout2774,
   input         cfg_dout2775,
   input         cfg_dout2776,
   input         cfg_dout2777,
   input         cfg_dout2778,
   input         cfg_dout2779,
   input         cfg_dout2780,
   input         cfg_dout2781,
   input         cfg_dout2782,
   input         cfg_dout2783,
   input         cfg_dout2784,
   input         cfg_dout2785,
   input         cfg_dout2786,
   input         cfg_dout2787,
   input         cfg_dout2788,
   input         cfg_dout2789,
   input         cfg_dout2790,
   input         cfg_dout2791,
   input         cfg_dout2792,
   input         cfg_dout2793,
   input         cfg_dout2794,
   input         cfg_dout2795,
   input         cfg_dout2796,
   input         cfg_dout2797,
   input         cfg_dout2798,
   input         cfg_dout2799,
   input         cfg_dout2800,
   input         cfg_dout2801,
   input         cfg_dout2802,
   input         cfg_dout2803,
   input         cfg_dout2804,
   input         cfg_dout2805,
   input         cfg_dout2806,
   input         cfg_dout2807,
   input         cfg_dout2808,
   input         cfg_dout2809,
   input         cfg_dout2810,
   input         cfg_dout2811,
   input         cfg_dout2812,
   input         cfg_dout2813,
   input         cfg_dout2814,
   input         cfg_dout2815,
   input         cfg_dout2816,
   input         cfg_dout2817,
   input         cfg_dout2818,
   input         cfg_dout2819,
   input         cfg_dout2820,
   input         cfg_dout2821,
   input         cfg_dout2822,
   input         cfg_dout2823,
   input         cfg_dout2824,
   input         cfg_dout2825,
   input         cfg_dout2826,
   input         cfg_dout2827,
   input         cfg_dout2828,
   input         cfg_dout2829,
   input         cfg_dout2830,
   input         cfg_dout2831,
   input         cfg_dout2832,
   input         cfg_dout2833,
   input         cfg_dout2834,
   input         cfg_dout2835,
   input         cfg_dout2836,
   input         cfg_dout2837,
   input         cfg_dout2838,
   input         cfg_dout2839,
   input         cfg_dout2840,
   input         cfg_dout2841,
   input         cfg_dout2842,
   input         cfg_dout2843,
   input         cfg_dout2844,
   input         cfg_dout2845,
   input         cfg_dout2846,
   input         cfg_dout2847,
   input         cfg_dout2848,
   input         cfg_dout2849,
   input         cfg_dout2850,
   input         cfg_dout2851,
   input         cfg_dout2852,
   input         cfg_dout2853,
   input         cfg_dout2854,
   input         cfg_dout2855,
   input         cfg_dout2856,
   input         cfg_dout2857,
   input         cfg_dout2858,
   input         cfg_dout2859,
   input         cfg_dout2860,
   input         cfg_dout2861,
   input         cfg_dout2862,
   input         cfg_dout2863,
   input         cfg_dout2864,
   input         cfg_dout2865,
   input         cfg_dout2866,
   input         cfg_dout2867,
   input         cfg_dout2868,
   input         cfg_dout2869,
   input         cfg_dout2870,
   input         cfg_dout2871,
   input         cfg_dout2872,
   input         cfg_dout2873,
   input         cfg_dout2874,
   input         cfg_dout2875,
   input         cfg_dout2876,
   input         cfg_dout2877,
   input         cfg_dout2878,
   input         cfg_dout2879,
   input         cfg_dout2880,
   input         cfg_dout2881,
   input         cfg_dout2882,
   input         cfg_dout2883,
   input         cfg_dout2884,
   input         cfg_dout2885,
   input         cfg_dout2886,
   input         cfg_dout2887,
   input         cfg_dout2888,
   input         cfg_dout2889,
   input         cfg_dout2890,
   input         cfg_dout2891,
   input         cfg_dout2892,
   input         cfg_dout2893,
   input         cfg_dout2894,
   input         cfg_dout2895,
   input         cfg_dout2896,
   input         cfg_dout2897,
   input         cfg_dout2898,
   input         cfg_dout2899,
   input         cfg_dout2900,
   input         cfg_dout2901,
   input         cfg_dout2902,
   input         cfg_dout2903,
   input         cfg_dout2904,
   input         cfg_dout2905,
   input         cfg_dout2906,
   input         cfg_dout2907,
   input         cfg_dout2908,
   input         cfg_dout2909,
   input         cfg_dout2910,
   input         cfg_dout2911,
   input         cfg_dout2912,
   input         cfg_dout2913,
   input         cfg_dout2914,
   input         cfg_dout2915,
   input         cfg_dout2916,
   input         cfg_dout2917,
   input         cfg_dout2918,
   input         cfg_dout2919,
   input         cfg_dout2920,
   input         cfg_dout2921,
   input         cfg_dout2922,
   input         cfg_dout2923,
   input         cfg_dout2924,
   input         cfg_dout2925,
   input         cfg_dout2926,
   input         cfg_dout2927,
   input         cfg_dout2928,
   input         cfg_dout2929,
   input         cfg_dout2930,
   input         cfg_dout2931,
   input         cfg_dout2932,
   input         cfg_dout2933,
   input         cfg_dout2934,
   input         cfg_dout2935,
   input         cfg_dout2936,
   input         cfg_dout2937,
   input         cfg_dout2938,
   input         cfg_dout2939,
   input         cfg_dout2940,
   input         cfg_dout2941,
   input         cfg_dout2942,
   input         cfg_dout2943,
   input         cfg_dout2944,
   input         cfg_dout2945,
   input         cfg_dout2946,
   input         cfg_dout2947,
   input         cfg_dout2948,
   input         cfg_dout2949,
   input         cfg_dout2950,
   input         cfg_dout2951,
   input         cfg_dout2952,
   input         cfg_dout2953,
   input         cfg_dout2954,
   input         cfg_dout2955,
   input         cfg_dout2956,
   input         cfg_dout2957,
   input         cfg_dout2958,
   input         cfg_dout2959,
   input         cfg_dout2960,
   input         cfg_dout2961,
   input         cfg_dout2962,
   input         cfg_dout2963,
   input         cfg_dout2964,
   input         cfg_dout2965,
   input         cfg_dout2966,
   input         cfg_dout2967,
   input         cfg_dout2968,
   input         cfg_dout2969,
   input         cfg_dout2970,
   input         cfg_dout2971,
   input         cfg_dout2972,
   input         cfg_dout2973,
   input         cfg_dout2974,
   input         cfg_dout2975,
   input         cfg_dout2976,
   input         cfg_dout2977,
   input         cfg_dout2978,
   input         cfg_dout2979,
   input         cfg_dout2980,
   input         cfg_dout2981,
   input         cfg_dout2982,
   input         cfg_dout2983,
   input         cfg_dout2984,
   input         cfg_dout2985,
   input         cfg_dout2986,
   input         cfg_dout2987,
   input         cfg_dout2988,
   input         cfg_dout2989,
   input         cfg_dout2990,
   input         cfg_dout2991,
   input         cfg_dout2992,
   input         cfg_dout2993,
   input         cfg_dout2994,
   input         cfg_dout2995,
   input         cfg_dout2996,
   input         cfg_dout2997,
   input         cfg_dout2998,
   input         cfg_dout2999,
   input         cfg_dout3000,
   input         cfg_dout3001,
   input         cfg_dout3002,
   input         cfg_dout3003,
   input         cfg_dout3004,
   input         cfg_dout3005,
   input         cfg_dout3006,
   input         cfg_dout3007,
   input         cfg_dout3008,
   input         cfg_dout3009,
   input         cfg_dout3010,
   input         cfg_dout3011,
   input         cfg_dout3012,
   input         cfg_dout3013,
   input         cfg_dout3014,
   input         cfg_dout3015,
   input         cfg_dout3016,
   input         cfg_dout3017,
   input         cfg_dout3018,
   input         cfg_dout3019,
   input         cfg_dout3020,
   input         cfg_dout3021,
   input         cfg_dout3022,
   input         cfg_dout3023,
   input         cfg_dout3024,
   input         cfg_dout3025,
   input         cfg_dout3026,
   input         cfg_dout3027,
   input         cfg_dout3028,
   input         cfg_dout3029,
   input         cfg_dout3030,
   input         cfg_dout3031,
   input         cfg_dout3032,
   input         cfg_dout3033,
   input         cfg_dout3034,
   input         cfg_dout3035,
   input         cfg_dout3036,
   input         cfg_dout3037,
   input         cfg_dout3038,
   input         cfg_dout3039,
   input         cfg_dout3040,
   input         cfg_dout3041,
   input         cfg_dout3042,
   input         cfg_dout3043,
   input         cfg_dout3044,
   input         cfg_dout3045,
   input         cfg_dout3046,
   input         cfg_dout3047,
   input         cfg_dout3048,
   input         cfg_dout3049,
   input         cfg_dout3050,
   input         cfg_dout3051,
   input         cfg_dout3052,
   input         cfg_dout3053,
   input         cfg_dout3054,
   input         cfg_dout3055,
   input         cfg_dout3056,
   input         cfg_dout3057,
   input         cfg_dout3058,
   input         cfg_dout3059,
   input         cfg_dout3060,
   input         cfg_dout3061,
   input         cfg_dout3062,
   input         cfg_dout3063,
   input         cfg_dout3064,
   input         cfg_dout3065,
   input         cfg_dout3066,
   input         cfg_dout3067,
   input         cfg_dout3068,
   input         cfg_dout3069,
   input         cfg_dout3070,
   input         cfg_dout3071,
   input         cfg_dout3072,
   input         cfg_dout3073,
   input         cfg_dout3074,
   input         cfg_dout3075,
   input         cfg_dout3076,
   input         cfg_dout3077,
   input         cfg_dout3078,
   input         cfg_dout3079,
   input         cfg_dout3080,
   input         cfg_dout3081,
   input         cfg_dout3082,
   input         cfg_dout3083,
   input         cfg_dout3084,
   input         cfg_dout3085,
   input         cfg_dout3086,
   input         cfg_dout3087,
   input         cfg_dout3088,
   input         cfg_dout3089,
   input         cfg_dout3090,
   input         cfg_dout3091,
   input         cfg_dout3092,
   input         cfg_dout3093,
   input         cfg_dout3094,
   input         cfg_dout3095,
   input         cfg_dout3096,
   input         cfg_dout3097,
   input         cfg_dout3098,
   input         cfg_dout3099,
   input         cfg_dout3100,
   input         cfg_dout3101,
   input         cfg_dout3102,
   input         cfg_dout3103,
   input         cfg_dout3104,
   input         cfg_dout3105,
   input         cfg_dout3106,
   input         cfg_dout3107,
   input         cfg_dout3108,
   input         cfg_dout3109,
   input         cfg_dout3110,
   input         cfg_dout3111,
   input         cfg_dout3112,
   input         cfg_dout3113,
   input         cfg_dout3114,
   input         cfg_dout3115,
   input         cfg_dout3116,
   input         cfg_dout3117,
   input         cfg_dout3118,
   input         cfg_dout3119,
   input         cfg_dout3120,
   input         cfg_dout3121,
   input         cfg_dout3122,
   input         cfg_dout3123,
   input         cfg_dout3124,
   input         cfg_dout3125,
   input         cfg_dout3126,
   input         cfg_dout3127,
   input         cfg_dout3128,
   input         cfg_dout3129,
   input         cfg_dout3130,
   input         cfg_dout3131,
   input         cfg_dout3132,
   input         cfg_dout3133,
   input         cfg_dout3134,
   input         cfg_dout3135,
   input         cfg_dout3136,
   input         cfg_dout3137,
   input         cfg_dout3138,
   input         cfg_dout3139,
   input         cfg_dout3140,
   input         cfg_dout3141,
   input         cfg_dout3142,
   input         cfg_dout3143,
   input         cfg_dout3144,
   input         cfg_dout3145,
   input         cfg_dout3146,
   input         cfg_dout3147,
   input         cfg_dout3148,
   input         cfg_dout3149,
   input         cfg_dout3150,
   input         cfg_dout3151,
   input         cfg_dout3152,
   input         cfg_dout3153,
   input         cfg_dout3154,
   input         cfg_dout3155,
   input         cfg_dout3156,
   input         cfg_dout3157,
   input         cfg_dout3158,
   input         cfg_dout3159,
   input         cfg_dout3160,
   input         cfg_dout3161,
   input         cfg_dout3162,
   input         cfg_dout3163,
   input         cfg_dout3164,
   input         cfg_dout3165,
   input         cfg_dout3166,
   input         cfg_dout3167,
   input         cfg_dout3168,
   input         cfg_dout3169,
   input         cfg_dout3170,
   input         cfg_dout3171,
   input         cfg_dout3172,
   input         cfg_dout3173,
   input         cfg_dout3174,
   input         cfg_dout3175,
   input         cfg_dout3176,
   input         cfg_dout3177,
   input         cfg_dout3178,
   input         cfg_dout3179,
   input         cfg_dout3180,
   input         cfg_dout3181,
   input         cfg_dout3182,
   input         cfg_dout3183,
   input         cfg_dout3184,
   input         cfg_dout3185,
   input         cfg_dout3186,
   input         cfg_dout3187,
   input         cfg_dout3188,
   input         cfg_dout3189,
   input         cfg_dout3190,
   input         cfg_dout3191,
   input         cfg_dout3192,
   input         cfg_dout3193,
   input         cfg_dout3194,
   input         cfg_dout3195,
   input         cfg_dout3196,
   input         cfg_dout3197,
   input         cfg_dout3198,
   input         cfg_dout3199,
   input         cfg_dout3200,
   input         cfg_dout3201,
   input         cfg_dout3202,
   input         cfg_dout3203,
   input         cfg_dout3204,
   input         cfg_dout3205,
   input         cfg_dout3206,
   input         cfg_dout3207,
   input         cfg_dout3208,
   input         cfg_dout3209,
   input         cfg_dout3210,
   input         cfg_dout3211,
   input         cfg_dout3212,
   input         cfg_dout3213,
   input         cfg_dout3214,
   input         cfg_dout3215,
   input         cfg_dout3216,
   input         cfg_dout3217,
   input         cfg_dout3218,
   input         cfg_dout3219,
   input         cfg_dout3220,
   input         cfg_dout3221,
   input         cfg_dout3222,
   input         cfg_dout3223,
   input         cfg_dout3224,
   input         cfg_dout3225,
   input         cfg_dout3226,
   input         cfg_dout3227,
   input         cfg_dout3228,
   input         cfg_dout3229,
   input         cfg_dout3230,
   input         cfg_dout3231,
   input         cfg_dout3232,
   input         cfg_dout3233,
   input         cfg_dout3234,
   input         cfg_dout3235,
   input         cfg_dout3236,
   input         cfg_dout3237,
   input         cfg_dout3238,
   input         cfg_dout3239,
   input         cfg_dout3240,
   input         cfg_dout3241,
   input         cfg_dout3242,
   input         cfg_dout3243,
   input         cfg_dout3244,
   input         cfg_dout3245,
   input         cfg_dout3246,
   input         cfg_dout3247,
   input         cfg_dout3248,
   input         cfg_dout3249,
   input         cfg_dout3250,
   input         cfg_dout3251,
   input         cfg_dout3252,
   input         cfg_dout3253,
   input         cfg_dout3254,
   input         cfg_dout3255,
   input         cfg_dout3256,
   input         cfg_dout3257,
   input         cfg_dout3258,
   input         cfg_dout3259,
   input         cfg_dout3260,
   input         cfg_dout3261,
   input         cfg_dout3262,
   input         cfg_dout3263,
   input         cfg_dout3264,
   input         cfg_dout3265,
   input         cfg_dout3266,
   input         cfg_dout3267,
   input         cfg_dout3268,
   input         cfg_dout3269,
   input         cfg_dout3270,
   input         cfg_dout3271,
   input         cfg_dout3272,
   input         cfg_dout3273,
   input         cfg_dout3274,
   input         cfg_dout3275,
   input         cfg_dout3276,
   input         cfg_dout3277,
   input         cfg_dout3278,
   input         cfg_dout3279,
   input         cfg_dout3280,
   input         cfg_dout3281,
   input         cfg_dout3282,
   input         cfg_dout3283,
   input         cfg_dout3284,
   input         cfg_dout3285,
   input         cfg_dout3286,
   input         cfg_dout3287,
   input         cfg_dout3288,
   input         cfg_dout3289,
   input         cfg_dout3290,
   input         cfg_dout3291,
   input         cfg_dout3292,
   input         cfg_dout3293,
   input         cfg_dout3294,
   input         cfg_dout3295,
   input         cfg_dout3296,
   input         cfg_dout3297,
   input         cfg_dout3298,
   input         cfg_dout3299,
   input         cfg_dout3300,
   input         cfg_dout3301,
   input         cfg_dout3302,
   input         cfg_dout3303,
   input         cfg_dout3304,
   input         cfg_dout3305,
   input         cfg_dout3306,
   input         cfg_dout3307,
   input         cfg_dout3308,
   input         cfg_dout3309,
   input         cfg_dout3310,
   input         cfg_dout3311,
   input         cfg_dout3312,
   input         cfg_dout3313,
   input         cfg_dout3314,
   input         cfg_dout3315,
   input         cfg_dout3316,
   input         cfg_dout3317,
   input         cfg_dout3318,
   input         cfg_dout3319,
   input         cfg_dout3320,
   input         cfg_dout3321,
   input         cfg_dout3322,
   input         cfg_dout3323,
   input         cfg_dout3324,
   input         cfg_dout3325,
   input         cfg_dout3326,
   input         cfg_dout3327,
   input         cfg_dout3328,
   input         cfg_dout3329,
   input         cfg_dout3330,
   input         cfg_dout3331,
   input         cfg_dout3332,
   input         cfg_dout3333,
   input         cfg_dout3334,
   input         cfg_dout3335,
   input         cfg_dout3336,
   input         cfg_dout3337,
   input         cfg_dout3338,
   input         cfg_dout3339,
   input         cfg_dout3340,
   input         cfg_dout3341,
   input         cfg_dout3342,
   input         cfg_dout3343,
   input         cfg_dout3344,
   input         cfg_dout3345,
   input         cfg_dout3346,
   input         cfg_dout3347,
   input         cfg_dout3348,
   input         cfg_dout3349,
   input         cfg_dout3350,
   input         cfg_dout3351,
   input         cfg_dout3352,
   input         cfg_dout3353,
   input         cfg_dout3354,
   input         cfg_dout3355,
   input         cfg_dout3356,
   input         cfg_dout3357,
   input         cfg_dout3358,
   input         cfg_dout3359,
   input         cfg_dout3360,
   input         cfg_dout3361,
   input         cfg_dout3362,
   input         cfg_dout3363,
   input         cfg_dout3364,
   input         cfg_dout3365,
   input         cfg_dout3366,
   input         cfg_dout3367,
   input         cfg_dout3368,
   input         cfg_dout3369,
   input         cfg_dout3370,
   input         cfg_dout3371,
   input         cfg_dout3372,
   input         cfg_dout3373,
   input         cfg_dout3374,
   input         cfg_dout3375,
   input         cfg_dout3376,
   input         cfg_dout3377,
   input         cfg_dout3378,
   input         cfg_dout3379,
   input         cfg_dout3380,
   input         cfg_dout3381,
   input         cfg_dout3382,
   input         cfg_dout3383,
   input         cfg_dout3384,
   input         cfg_dout3385,
   input         cfg_dout3386,
   input         cfg_dout3387,
   input         cfg_dout3388,
   input         cfg_dout3389,
   input         cfg_dout3390,
   input         cfg_dout3391,
   input         cfg_dout3392,
   input         cfg_dout3393,
   input         cfg_dout3394,
   input         cfg_dout3395,
   input         cfg_dout3396,
   input         cfg_dout3397,
   input         cfg_dout3398,
   input         cfg_dout3399,
   input         cfg_dout3400,
   input         cfg_dout3401,
   input         cfg_dout3402,
   input         cfg_dout3403,
   input         cfg_dout3404,
   input         cfg_dout3405,
   input         cfg_dout3406,
   input         cfg_dout3407,
   input         cfg_dout3408,
   input         cfg_dout3409,
   input         cfg_dout3410,
   input         cfg_dout3411,
   input         cfg_dout3412,
   input         cfg_dout3413,
   input         cfg_dout3414,
   input         cfg_dout3415,
   input         cfg_dout3416,
   input         cfg_dout3417,
   input         cfg_dout3418,
   input         cfg_dout3419,
   input         cfg_dout3420,
   input         cfg_dout3421,
   input         cfg_dout3422,
   input         cfg_dout3423,
   input         cfg_dout3424,
   input         cfg_dout3425,
   input         cfg_dout3426,
   input         cfg_dout3427,
   input         cfg_dout3428,
   input         cfg_dout3429,
   input         cfg_dout3430,
   input         cfg_dout3431,
   input         cfg_dout3432,
   input         cfg_dout3433,
   input         cfg_dout3434,
   input         cfg_dout3435,
   input         cfg_dout3436,
   input         cfg_dout3437,
   input         cfg_dout3438,
   input         cfg_dout3439,
   input         cfg_dout3440,
   input         cfg_dout3441,
   input         cfg_dout3442,
   input         cfg_dout3443,
   input         cfg_dout3444,
   input         cfg_dout3445,
   input         cfg_dout3446,
   input         cfg_dout3447,
   input         cfg_dout3448,
   input         cfg_dout3449,
   input         cfg_dout3450,
   input         cfg_dout3451,
   input         cfg_dout3452,
   input         cfg_dout3453,
   input         cfg_dout3454,
   input         cfg_dout3455,
   input         cfg_dout3456,
   input         cfg_dout3457,
   input         cfg_dout3458,
   input         cfg_dout3459,
   input         cfg_dout3460,
   input         cfg_dout3461,
   input         cfg_dout3462,
   input         cfg_dout3463,
   input         cfg_dout3464,
   input         cfg_dout3465,
   input         cfg_dout3466,
   input         cfg_dout3467,
   input         cfg_dout3468,
   input         cfg_dout3469,
   input         cfg_dout3470,
   input         cfg_dout3471,
   input         cfg_dout3472,
   input         cfg_dout3473,
   input         cfg_dout3474,
   input         cfg_dout3475,
   input         cfg_dout3476,
   input         cfg_dout3477,
   input         cfg_dout3478,
   input         cfg_dout3479,
   input         cfg_dout3480,
   input         cfg_dout3481,
   input         cfg_dout3482,
   input         cfg_dout3483,
   input         cfg_dout3484,
   input         cfg_dout3485,
   input         cfg_dout3486,
   input         cfg_dout3487,
   input         cfg_dout3488,
   input         cfg_dout3489,
   input         cfg_dout3490,
   input         cfg_dout3491,
   input         cfg_dout3492,
   input         cfg_dout3493,
   input         cfg_dout3494,
   input         cfg_dout3495,
   input         cfg_dout3496,
   input         cfg_dout3497,
   input         cfg_dout3498,
   input         cfg_dout3499,
   input         cfg_dout3500,
   input         cfg_dout3501,
   input         cfg_dout3502,
   input         cfg_dout3503,
   input         cfg_dout3504,
   input         cfg_dout3505,
   input         cfg_dout3506,
   input         cfg_dout3507,
   input         cfg_dout3508,
   input         cfg_dout3509,
   input         cfg_dout3510,
   input         cfg_dout3511,
   input         cfg_dout3512,
   input         cfg_dout3513,
   input         cfg_dout3514,
   input         cfg_dout3515,
   input         cfg_dout3516,
   input         cfg_dout3517,
   input         cfg_dout3518,
   input         cfg_dout3519,
   input         cfg_dout3520,
   input         cfg_dout3521,
   input         cfg_dout3522,
   input         cfg_dout3523,
   input         cfg_dout3524,
   input         cfg_dout3525,
   input         cfg_dout3526,
   input         cfg_dout3527,
   input         cfg_dout3528,
   input         cfg_dout3529,
   input         cfg_dout3530,
   input         cfg_dout3531,
   input         cfg_dout3532,
   input         cfg_dout3533,
   input         cfg_dout3534,
   input         cfg_dout3535,
   input         cfg_dout3536,
   input         cfg_dout3537,
   input         cfg_dout3538,
   input         cfg_dout3539,
   input         cfg_dout3540,
   input         cfg_dout3541,
   input         cfg_dout3542,
   input         cfg_dout3543,
   input         cfg_dout3544,
   input         cfg_dout3545,
   input         cfg_dout3546,
   input         cfg_dout3547,
   input         cfg_dout3548,
   input         cfg_dout3549,
   input         cfg_dout3550,
   input         cfg_dout3551,
   input         cfg_dout3552,
   input         cfg_dout3553,
   input         cfg_dout3554,
   input         cfg_dout3555,
   input         cfg_dout3556,
   input         cfg_dout3557,
   input         cfg_dout3558,
   input         cfg_dout3559,
   input         cfg_dout3560,
   input         cfg_dout3561,
   input         cfg_dout3562,
   input         cfg_dout3563,
   input         cfg_dout3564,
   input         cfg_dout3565,
   input         cfg_dout3566,
   input         cfg_dout3567,
   input         cfg_dout3568,
   input         cfg_dout3569,
   input         cfg_dout3570,
   input         cfg_dout3571,
   input         cfg_dout3572,
   input         cfg_dout3573,
   input         cfg_dout3574,
   input         cfg_dout3575,
   input         cfg_dout3576,
   input         cfg_dout3577,
   input         cfg_dout3578,
   input         cfg_dout3579,
   input         cfg_dout3580,
   input         cfg_dout3581,
   input         cfg_dout3582,
   input         cfg_dout3583,
   input         cfg_dout3584,
   input         cfg_dout3585,
   input         cfg_dout3586,
   input         cfg_dout3587,
   input         cfg_dout3588,
   input         cfg_dout3589,
   input         cfg_dout3590,
   input         cfg_dout3591,
   input         cfg_dout3592,
   input         cfg_dout3593,
   input         cfg_dout3594,
   input         cfg_dout3595,
   input         cfg_dout3596,
   input         cfg_dout3597,
   input         cfg_dout3598,
   input         cfg_dout3599,
   input         cfg_dout3600,
   input         cfg_dout3601,
   input         cfg_dout3602,
   input         cfg_dout3603,
   input         cfg_dout3604,
   input         cfg_dout3605,
   input         cfg_dout3606,
   input         cfg_dout3607,
   input         cfg_dout3608,
   input         cfg_dout3609,
   input         cfg_dout3610,
   input         cfg_dout3611,
   input         cfg_dout3612,
   input         cfg_dout3613,
   input         cfg_dout3614,
   input         cfg_dout3615,
   input         cfg_dout3616,
   input         cfg_dout3617,
   input         cfg_dout3618,
   input         cfg_dout3619,
   input         cfg_dout3620,
   input         cfg_dout3621,
   input         cfg_dout3622,
   input         cfg_dout3623,
   input         cfg_dout3624,
   input         cfg_dout3625,
   input         cfg_dout3626,
   input         cfg_dout3627,
   input         cfg_dout3628,
   input         cfg_dout3629,
   input         cfg_dout3630,
   input         cfg_dout3631,
   input         cfg_dout3632,
   input         cfg_dout3633,
   input         cfg_dout3634,
   input         cfg_dout3635,
   input         cfg_dout3636,
   input         cfg_dout3637,
   input         cfg_dout3638,
   input         cfg_dout3639,
   input         cfg_dout3640,
   input         cfg_dout3641,
   input         cfg_dout3642,
   input         cfg_dout3643,
   input         cfg_dout3644,
   input         cfg_dout3645,
   input         cfg_dout3646,
   input         cfg_dout3647,
   input         cfg_dout3648,
   input         cfg_dout3649,
   input         cfg_dout3650,
   input         cfg_dout3651,
   input         cfg_dout3652,
   input         cfg_dout3653,
   input         cfg_dout3654,
   input         cfg_dout3655,
   input         cfg_dout3656,
   input         cfg_dout3657,
   input         cfg_dout3658,
   input         cfg_dout3659,
   input         cfg_dout3660,
   input         cfg_dout3661,
   input         cfg_dout3662,
   input         cfg_dout3663,
   input         cfg_dout3664,
   input         cfg_dout3665,
   input         cfg_dout3666,
   input         cfg_dout3667,
   input         cfg_dout3668,
   input         cfg_dout3669,
   input         cfg_dout3670,
   input         cfg_dout3671,
   input         cfg_dout3672,
   input         cfg_dout3673,
   input         cfg_dout3674,
   input         cfg_dout3675,
   input         cfg_dout3676,
   input         cfg_dout3677,
   input         cfg_dout3678,
   input         cfg_dout3679,
   input         cfg_dout3680,
   input         cfg_dout3681,
   input         cfg_dout3682,
   input         cfg_dout3683,
   input         cfg_dout3684,
   input         cfg_dout3685,
   input         cfg_dout3686,
   input         cfg_dout3687,
   input         cfg_dout3688,
   input         cfg_dout3689,
   input         cfg_dout3690,
   input         cfg_dout3691,
   input         cfg_dout3692,
   input         cfg_dout3693,
   input         cfg_dout3694,
   input         cfg_dout3695,
   input         cfg_dout3696,
   input         cfg_dout3697,
   input         cfg_dout3698,
   input         cfg_dout3699,
   input         cfg_dout3700,
   input         cfg_dout3701,
   input         cfg_dout3702,
   input         cfg_dout3703,
   input         cfg_dout3704,
   input         cfg_dout3705,
   input         cfg_dout3706,
   input         cfg_dout3707,
   input         cfg_dout3708,
   input         cfg_dout3709,
   input         cfg_dout3710,
   input         cfg_dout3711,
   input         cfg_dout3712,
   input         cfg_dout3713,
   input         cfg_dout3714,
   input         cfg_dout3715,
   input         cfg_dout3716,
   input         cfg_dout3717,
   input         cfg_dout3718,
   input         cfg_dout3719,
   input         cfg_dout3720,
   input         cfg_dout3721,
   input         cfg_dout3722,
   input         cfg_dout3723,
   input         cfg_dout3724,
   input         cfg_dout3725,
   input         cfg_dout3726,
   input         cfg_dout3727,
   input         cfg_dout3728,
   input         cfg_dout3729,
   input         cfg_dout3730,
   input         cfg_dout3731,
   input         cfg_dout3732,
   input         cfg_dout3733,
   input         cfg_dout3734,
   input         cfg_dout3735,
   input         cfg_dout3736,
   input         cfg_dout3737,
   input         cfg_dout3738,
   input         cfg_dout3739,
   input         cfg_dout3740,
   input         cfg_dout3741,
   input         cfg_dout3742,
   input         cfg_dout3743,
   input         cfg_dout3744,
   input         cfg_dout3745,
   input         cfg_dout3746,
   input         cfg_dout3747,
   input         cfg_dout3748,
   input         cfg_dout3749,
   input         cfg_dout3750,
   input         cfg_dout3751,
   input         cfg_dout3752,
   input         cfg_dout3753,
   input         cfg_dout3754,
   input         cfg_dout3755,
   input         cfg_dout3756,
   input         cfg_dout3757,
   input         cfg_dout3758,
   input         cfg_dout3759,
   input         cfg_dout3760,
   input         cfg_dout3761,
   input         cfg_dout3762,
   input         cfg_dout3763,
   input         cfg_dout3764,
   input         cfg_dout3765,
   input         cfg_dout3766,
   input         cfg_dout3767,
   input         cfg_dout3768,
   input         cfg_dout3769,
   input         cfg_dout3770,
   input         cfg_dout3771,
   input         cfg_dout3772,
   input         cfg_dout3773,
   input         cfg_dout3774,
   input         cfg_dout3775,
   input         cfg_dout3776,
   input         cfg_dout3777,
   input         cfg_dout3778,
   input         cfg_dout3779,
   input         cfg_dout3780,
   input         cfg_dout3781,
   input         cfg_dout3782,
   input         cfg_dout3783,
   input         cfg_dout3784,
   input         cfg_dout3785,
   input         cfg_dout3786,
   input         cfg_dout3787,
   input         cfg_dout3788,
   input         cfg_dout3789,
   input         cfg_dout3790,
   input         cfg_dout3791,
   input         cfg_dout3792,
   input         cfg_dout3793,
   input         cfg_dout3794,
   input         cfg_dout3795,
   input         cfg_dout3796,
   input         cfg_dout3797,
   input         cfg_dout3798,
   input         cfg_dout3799,
   input         cfg_dout3800,
   input         cfg_dout3801,
   input         cfg_dout3802,
   input         cfg_dout3803,
   input         cfg_dout3804,
   input         cfg_dout3805,
   input         cfg_dout3806,
   input         cfg_dout3807,
   input         cfg_dout3808,
   input         cfg_dout3809,
   input         cfg_dout3810,
   input         cfg_dout3811,
   input         cfg_dout3812,
   input         cfg_dout3813,
   input         cfg_dout3814,
   input         cfg_dout3815,
   input         cfg_dout3816,
   input         cfg_dout3817,
   input         cfg_dout3818,
   input         cfg_dout3819,
   input         cfg_dout3820,
   input         cfg_dout3821,
   input         cfg_dout3822,
   input         cfg_dout3823,
   input         cfg_dout3824,
   input         cfg_dout3825,
   input         cfg_dout3826,
   input         cfg_dout3827,
   input         cfg_dout3828,
   input         cfg_dout3829,
   input         cfg_dout3830,
   input         cfg_dout3831,
   input         cfg_dout3832,
   input         cfg_dout3833,
   input         cfg_dout3834,
   input         cfg_dout3835,
   input         cfg_dout3836,
   input         cfg_dout3837,
   input         cfg_dout3838,
   input         cfg_dout3839,
   input         cfg_dout3840,
   input         cfg_dout3841,
   input         cfg_dout3842,
   input         cfg_dout3843,
   input         cfg_dout3844,
   input         cfg_dout3845,
   input         cfg_dout3846,
   input         cfg_dout3847,
   input         cfg_dout3848,
   input         cfg_dout3849,
   input         cfg_dout3850,
   input         cfg_dout3851,
   input         cfg_dout3852,
   input         cfg_dout3853,
   input         cfg_dout3854,
   input         cfg_dout3855,
   input         cfg_dout3856,
   input         cfg_dout3857,
   input         cfg_dout3858,
   input         cfg_dout3859,
   input         cfg_dout3860,
   input         cfg_dout3861,
   input         cfg_dout3862,
   input         cfg_dout3863,
   input         cfg_dout3864,
   input         cfg_dout3865,
   input         cfg_dout3866,
   input         cfg_dout3867,
   input         cfg_dout3868,
   input         cfg_dout3869,
   input         cfg_dout3870,
   input         cfg_dout3871,
   input         cfg_dout3872,
   input         cfg_dout3873,
   input         cfg_dout3874,
   input         cfg_dout3875,
   input         cfg_dout3876,
   input         cfg_dout3877,
   input         cfg_dout3878,
   input         cfg_dout3879,
   input         cfg_dout3880,
   input         cfg_dout3881,
   input         cfg_dout3882,
   input         cfg_dout3883,
   input         cfg_dout3884,
   input         cfg_dout3885,
   input         cfg_dout3886,
   input         cfg_dout3887,
   input         cfg_dout3888,
   input         cfg_dout3889,
   input         cfg_dout3890,
   input         cfg_dout3891,
   input         cfg_dout3892,
   input         cfg_dout3893,
   input         cfg_dout3894,
   input         cfg_dout3895,
   input         cfg_dout3896,
   input         cfg_dout3897,
   input         cfg_dout3898,
   input         cfg_dout3899,
   input         cfg_dout3900,
   input         cfg_dout3901,
   input         cfg_dout3902,
   input         cfg_dout3903,
   input         cfg_dout3904,
   input         cfg_dout3905,
   input         cfg_dout3906,
   input         cfg_dout3907,
   input         cfg_dout3908,
   input         cfg_dout3909,
   input         cfg_dout3910,
   input         cfg_dout3911,
   input         cfg_dout3912,
   input         cfg_dout3913,
   input         cfg_dout3914,
   input         cfg_dout3915,
   input         cfg_dout3916,
   input         cfg_dout3917,
   input         cfg_dout3918,
   input         cfg_dout3919,
   input         cfg_dout3920,
   input         cfg_dout3921,
   input         cfg_dout3922,
   input         cfg_dout3923,
   input         cfg_dout3924,
   input         cfg_dout3925,
   input         cfg_dout3926,
   input         cfg_dout3927,
   input         cfg_dout3928,
   input         cfg_dout3929,
   input         cfg_dout3930,
   input         cfg_dout3931,
   input         cfg_dout3932,
   input         cfg_dout3933,
   input         cfg_dout3934,
   input         cfg_dout3935,
   input         cfg_dout3936,
   input         cfg_dout3937,
   input         cfg_dout3938,
   input         cfg_dout3939,
   input         cfg_dout3940,
   input         cfg_dout3941,
   input         cfg_dout3942,
   input         cfg_dout3943,
   input         cfg_dout3944,
   input         cfg_dout3945,
   input         cfg_dout3946,
   input         cfg_dout3947,
   input         cfg_dout3948,
   input         cfg_dout3949,
   input         cfg_dout3950,
   input         cfg_dout3951,
   input         cfg_dout3952,
   input         cfg_dout3953,
   input         cfg_dout3954,
   input         cfg_dout3955,
   input         cfg_dout3956,
   input         cfg_dout3957,
   input         cfg_dout3958,
   input         cfg_dout3959,
   input         cfg_dout3960,
   input         cfg_dout3961,
   input         cfg_dout3962,
   input         cfg_dout3963,
   input         cfg_dout3964,
   input         cfg_dout3965,
   input         cfg_dout3966,
   input         cfg_dout3967,
   input         cfg_dout3968,
   input         cfg_dout3969,
   input         cfg_dout3970,
   input         cfg_dout3971,
   input         cfg_dout3972,
   input         cfg_dout3973,
   input         cfg_dout3974,
   input         cfg_dout3975,
   input         cfg_dout3976,
   input         cfg_dout3977,
   input         cfg_dout3978,
   input         cfg_dout3979,
   input         cfg_dout3980,
   input         cfg_dout3981,
   input         cfg_dout3982,
   input         cfg_dout3983,
   input         cfg_dout3984,
   input         cfg_dout3985,
   input         cfg_dout3986,
   input         cfg_dout3987,
   input         cfg_dout3988,
   input         cfg_dout3989,
   input         cfg_dout3990,
   input         cfg_dout3991,
   input         cfg_dout3992,
   input         cfg_dout3993,
   input         cfg_dout3994,
   input         cfg_dout3995,
   input         cfg_dout3996,
   input         cfg_dout3997,
   input         cfg_dout3998,
   input         cfg_dout3999,
   input         cfg_dout4000,
   input         cfg_dout4001,
   input         cfg_dout4002,
   input         cfg_dout4003,
   input         cfg_dout4004,
   input         cfg_dout4005,
   input         cfg_dout4006,
   input         cfg_dout4007,
   input         cfg_dout4008,
   input         cfg_dout4009,
   input         cfg_dout4010,
   input         cfg_dout4011,
   input         cfg_dout4012,
   input         cfg_dout4013,
   input         cfg_dout4014,
   input         cfg_dout4015,
   input         cfg_dout4016,
   input         cfg_dout4017,
   input         cfg_dout4018,
   input         cfg_dout4019,
   input         cfg_dout4020,
   input         cfg_dout4021,
   input         cfg_dout4022,
   input         cfg_dout4023,
   input         cfg_dout4024,
   input         cfg_dout4025,
   input         cfg_dout4026,
   input         cfg_dout4027,
   input         cfg_dout4028,
   input         cfg_dout4029,
   input         cfg_dout4030,
   input         cfg_dout4031,
   input         cfg_dout4032,
   input         cfg_dout4033,
   input         cfg_dout4034,
   input         cfg_dout4035,
   input         cfg_dout4036,
   input         cfg_dout4037,
   input         cfg_dout4038,
   input         cfg_dout4039,
   input         cfg_dout4040,
   input         cfg_dout4041,
   input         cfg_dout4042,
   input         cfg_dout4043,
   input         cfg_dout4044,
   input         cfg_dout4045,
   input         cfg_dout4046,
   input         cfg_dout4047,
   input         cfg_dout4048,
   input         cfg_dout4049,
   input         cfg_dout4050,
   input         cfg_dout4051,
   input         cfg_dout4052,
   input         cfg_dout4053,
   input         cfg_dout4054,
   input         cfg_dout4055,
   input         cfg_dout4056,
   input         cfg_dout4057,
   input         cfg_dout4058,
   input         cfg_dout4059,
   input         cfg_dout4060,
   input         cfg_dout4061,
   input         cfg_dout4062,
   input         cfg_dout4063,
   input         cfg_dout4064,
   input         cfg_dout4065,
   input         cfg_dout4066,
   input         cfg_dout4067,
   input         cfg_dout4068,
   input         cfg_dout4069,
   input         cfg_dout4070,
   input         cfg_dout4071,
   input         cfg_dout4072,
   input         cfg_dout4073,
   input         cfg_dout4074,
   input         cfg_dout4075,
   input         cfg_dout4076,
   input         cfg_dout4077,
   input         cfg_dout4078,
   input         cfg_dout4079,
   input         cfg_dout4080,
   input         cfg_dout4081,
   input         cfg_dout4082,
   input         cfg_dout4083,
   input         cfg_dout4084,
   input         cfg_dout4085,
   input         cfg_dout4086,
   input         cfg_dout4087,
   input         cfg_dout4088,
   input         cfg_dout4089,
   input         cfg_dout4090,
   input         cfg_dout4091,
   input         cfg_dout4092,
   input         cfg_dout4093,
   input         cfg_dout4094,
   input         cfg_dout4095,
   input         tc_cfg_dout,
   input         cc_cfg_dout0,
   input         cc_cfg_dout1,
   input         cc_cfg_dout2,
   input         cc_cfg_dout3,
   input         match_out0,
   input         match_out1,
   input         match_out2,
   input         match_out3,
   input         match_out4,
   input         match_out5,
   input         match_out6,
   input         match_out7,
   input         match_out8,
   input         match_out9,
   input         match_out10,
   input         match_out11,
   input         match_out12,
   input         match_out13,
   input         match_out14,
   input         match_out15,
   input         match_out16,
   input         match_out17,
   input         match_out18,
   input         match_out19,
   input         match_out20,
   input         match_out21,
   input         match_out22,
   input         match_out23,
   input         match_out24,
   input         match_out25,
   input         match_out26,
   input         match_out27,
   input         match_out28,
   input         match_out29,
   input         match_out30,
   input         match_out31,
   input         match_out32,
   input         match_out33,
   input         match_out34,
   input         match_out35,
   input         match_out36,
   input         match_out37,
   input         match_out38,
   input         match_out39,
   input         match_out40,
   input         match_out41,
   input         match_out42,
   input         match_out43,
   input         match_out44,
   input         match_out45,
   input         match_out46,
   input         match_out47,
   input         match_out48,
   input         match_out49,
   input         match_out50,
   input         match_out51,
   input         match_out52,
   input         match_out53,
   input         match_out54,
   input         match_out55,
   input         match_out56,
   input         match_out57,
   input         match_out58,
   input         match_out59,
   input         match_out60,
   input         match_out61,
   input         match_out62,
   input         match_out63,
   input         match_out64,
   input         match_out65,
   input         match_out66,
   input         match_out67,
   input         match_out68,
   input         match_out69,
   input         match_out70,
   input         match_out71,
   input         match_out72,
   input         match_out73,
   input         match_out74,
   input         match_out75,
   input         match_out76,
   input         match_out77,
   input         match_out78,
   input         match_out79,
   input         match_out80,
   input         match_out81,
   input         match_out82,
   input         match_out83,
   input         match_out84,
   input         match_out85,
   input         match_out86,
   input         match_out87,
   input         match_out88,
   input         match_out89,
   input         match_out90,
   input         match_out91,
   input         match_out92,
   input         match_out93,
   input         match_out94,
   input         match_out95,
   input         match_out96,
   input         match_out97,
   input         match_out98,
   input         match_out99,
   input         match_out100,
   input         match_out101,
   input         match_out102,
   input         match_out103,
   input         match_out104,
   input         match_out105,
   input         match_out106,
   input         match_out107,
   input         match_out108,
   input         match_out109,
   input         match_out110,
   input         match_out111,
   input         match_out112,
   input         match_out113,
   input         match_out114,
   input         match_out115,
   input         match_out116,
   input         match_out117,
   input         match_out118,
   input         match_out119,
   input         match_out120,
   input         match_out121,
   input         match_out122,
   input         match_out123,
   input         match_out124,
   input         match_out125,
   input         match_out126,
   input         match_out127,
   input         match_out128,
   input         match_out129,
   input         match_out130,
   input         match_out131,
   input         match_out132,
   input         match_out133,
   input         match_out134,
   input         match_out135,
   input         match_out136,
   input         match_out137,
   input         match_out138,
   input         match_out139,
   input         match_out140,
   input         match_out141,
   input         match_out142,
   input         match_out143,
   input         match_out144,
   input         match_out145,
   input         match_out146,
   input         match_out147,
   input         match_out148,
   input         match_out149,
   input         match_out150,
   input         match_out151,
   input         match_out152,
   input         match_out153,
   input         match_out154,
   input         match_out155,
   input         match_out156,
   input         match_out157,
   input         match_out158,
   input         match_out159,
   input         match_out160,
   input         match_out161,
   input         match_out162,
   input         match_out163,
   input         match_out164,
   input         match_out165,
   input         match_out166,
   input         match_out167,
   input         match_out168,
   input         match_out169,
   input         match_out170,
   input         match_out171,
   input         match_out172,
   input         match_out173,
   input         match_out174,
   input         match_out175,
   input         match_out176,
   input         match_out177,
   input         match_out178,
   input         match_out179,
   input         match_out180,
   input         match_out181,
   input         match_out182,
   input         match_out183,
   input         match_out184,
   input         match_out185,
   input         match_out186,
   input         match_out187,
   input         match_out188,
   input         match_out189,
   input         match_out190,
   input         match_out191,
   input         match_out192,
   input         match_out193,
   input         match_out194,
   input         match_out195,
   input         match_out196,
   input         match_out197,
   input         match_out198,
   input         match_out199,
   input         match_out200,
   input         match_out201,
   input         match_out202,
   input         match_out203,
   input         match_out204,
   input         match_out205,
   input         match_out206,
   input         match_out207,
   input         match_out208,
   input         match_out209,
   input         match_out210,
   input         match_out211,
   input         match_out212,
   input         match_out213,
   input         match_out214,
   input         match_out215,
   input         match_out216,
   input         match_out217,
   input         match_out218,
   input         match_out219,
   input         match_out220,
   input         match_out221,
   input         match_out222,
   input         match_out223,
   input         match_out224,
   input         match_out225,
   input         match_out226,
   input         match_out227,
   input         match_out228,
   input         match_out229,
   input         match_out230,
   input         match_out231,
   input         match_out232,
   input         match_out233,
   input         match_out234,
   input         match_out235,
   input         match_out236,
   input         match_out237,
   input         match_out238,
   input         match_out239,
   input         match_out240,
   input         match_out241,
   input         match_out242,
   input         match_out243,
   input         match_out244,
   input         match_out245,
   input         match_out246,
   input         match_out247,
   input         match_out248,
   input         match_out249,
   input         match_out250,
   input         match_out251,
   input         match_out252,
   input         match_out253,
   input         match_out254,
   input         match_out255,
   input         match_out256,
   input         match_out257,
   input         match_out258,
   input         match_out259,
   input         match_out260,
   input         match_out261,
   input         match_out262,
   input         match_out263,
   input         match_out264,
   input         match_out265,
   input         match_out266,
   input         match_out267,
   input         match_out268,
   input         match_out269,
   input         match_out270,
   input         match_out271,
   input         match_out272,
   input         match_out273,
   input         match_out274,
   input         match_out275,
   input         match_out276,
   input         match_out277,
   input         match_out278,
   input         match_out279,
   input         match_out280,
   input         match_out281,
   input         match_out282,
   input         match_out283,
   input         match_out284,
   input         match_out285,
   input         match_out286,
   input         match_out287,
   input         match_out288,
   input         match_out289,
   input         match_out290,
   input         match_out291,
   input         match_out292,
   input         match_out293,
   input         match_out294,
   input         match_out295,
   input         match_out296,
   input         match_out297,
   input         match_out298,
   input         match_out299,
   input         match_out300,
   input         match_out301,
   input         match_out302,
   input         match_out303,
   input         match_out304,
   input         match_out305,
   input         match_out306,
   input         match_out307,
   input         match_out308,
   input         match_out309,
   input         match_out310,
   input         match_out311,
   input         match_out312,
   input         match_out313,
   input         match_out314,
   input         match_out315,
   input         match_out316,
   input         match_out317,
   input         match_out318,
   input         match_out319,
   input         match_out320,
   input         match_out321,
   input         match_out322,
   input         match_out323,
   input         match_out324,
   input         match_out325,
   input         match_out326,
   input         match_out327,
   input         match_out328,
   input         match_out329,
   input         match_out330,
   input         match_out331,
   input         match_out332,
   input         match_out333,
   input         match_out334,
   input         match_out335,
   input         match_out336,
   input         match_out337,
   input         match_out338,
   input         match_out339,
   input         match_out340,
   input         match_out341,
   input         match_out342,
   input         match_out343,
   input         match_out344,
   input         match_out345,
   input         match_out346,
   input         match_out347,
   input         match_out348,
   input         match_out349,
   input         match_out350,
   input         match_out351,
   input         match_out352,
   input         match_out353,
   input         match_out354,
   input         match_out355,
   input         match_out356,
   input         match_out357,
   input         match_out358,
   input         match_out359,
   input         match_out360,
   input         match_out361,
   input         match_out362,
   input         match_out363,
   input         match_out364,
   input         match_out365,
   input         match_out366,
   input         match_out367,
   input         match_out368,
   input         match_out369,
   input         match_out370,
   input         match_out371,
   input         match_out372,
   input         match_out373,
   input         match_out374,
   input         match_out375,
   input         match_out376,
   input         match_out377,
   input         match_out378,
   input         match_out379,
   input         match_out380,
   input         match_out381,
   input         match_out382,
   input         match_out383,
   input         match_out384,
   input         match_out385,
   input         match_out386,
   input         match_out387,
   input         match_out388,
   input         match_out389,
   input         match_out390,
   input         match_out391,
   input         match_out392,
   input         match_out393,
   input         match_out394,
   input         match_out395,
   input         match_out396,
   input         match_out397,
   input         match_out398,
   input         match_out399,
   input         match_out400,
   input         match_out401,
   input         match_out402,
   input         match_out403,
   input         match_out404,
   input         match_out405,
   input         match_out406,
   input         match_out407,
   input         match_out408,
   input         match_out409,
   input         match_out410,
   input         match_out411,
   input         match_out412,
   input         match_out413,
   input         match_out414,
   input         match_out415,
   input         match_out416,
   input         match_out417,
   input         match_out418,
   input         match_out419,
   input         match_out420,
   input         match_out421,
   input         match_out422,
   input         match_out423,
   input         match_out424,
   input         match_out425,
   input         match_out426,
   input         match_out427,
   input         match_out428,
   input         match_out429,
   input         match_out430,
   input         match_out431,
   input         match_out432,
   input         match_out433,
   input         match_out434,
   input         match_out435,
   input         match_out436,
   input         match_out437,
   input         match_out438,
   input         match_out439,
   input         match_out440,
   input         match_out441,
   input         match_out442,
   input         match_out443,
   input         match_out444,
   input         match_out445,
   input         match_out446,
   input         match_out447,
   input         match_out448,
   input         match_out449,
   input         match_out450,
   input         match_out451,
   input         match_out452,
   input         match_out453,
   input         match_out454,
   input         match_out455,
   input         match_out456,
   input         match_out457,
   input         match_out458,
   input         match_out459,
   input         match_out460,
   input         match_out461,
   input         match_out462,
   input         match_out463,
   input         match_out464,
   input         match_out465,
   input         match_out466,
   input         match_out467,
   input         match_out468,
   input         match_out469,
   input         match_out470,
   input         match_out471,
   input         match_out472,
   input         match_out473,
   input         match_out474,
   input         match_out475,
   input         match_out476,
   input         match_out477,
   input         match_out478,
   input         match_out479,
   input         match_out480,
   input         match_out481,
   input         match_out482,
   input         match_out483,
   input         match_out484,
   input         match_out485,
   input         match_out486,
   input         match_out487,
   input         match_out488,
   input         match_out489,
   input         match_out490,
   input         match_out491,
   input         match_out492,
   input         match_out493,
   input         match_out494,
   input         match_out495,
   input         match_out496,
   input         match_out497,
   input         match_out498,
   input         match_out499,
   input         match_out500,
   input         match_out501,
   input         match_out502,
   input         match_out503,
   input         match_out504,
   input         match_out505,
   input         match_out506,
   input         match_out507,
   input         match_out508,
   input         match_out509,
   input         match_out510,
   input         match_out511,
   input         match_out512,
   input         match_out513,
   input         match_out514,
   input         match_out515,
   input         match_out516,
   input         match_out517,
   input         match_out518,
   input         match_out519,
   input         match_out520,
   input         match_out521,
   input         match_out522,
   input         match_out523,
   input         match_out524,
   input         match_out525,
   input         match_out526,
   input         match_out527,
   input         match_out528,
   input         match_out529,
   input         match_out530,
   input         match_out531,
   input         match_out532,
   input         match_out533,
   input         match_out534,
   input         match_out535,
   input         match_out536,
   input         match_out537,
   input         match_out538,
   input         match_out539,
   input         match_out540,
   input         match_out541,
   input         match_out542,
   input         match_out543,
   input         match_out544,
   input         match_out545,
   input         match_out546,
   input         match_out547,
   input         match_out548,
   input         match_out549,
   input         match_out550,
   input         match_out551,
   input         match_out552,
   input         match_out553,
   input         match_out554,
   input         match_out555,
   input         match_out556,
   input         match_out557,
   input         match_out558,
   input         match_out559,
   input         match_out560,
   input         match_out561,
   input         match_out562,
   input         match_out563,
   input         match_out564,
   input         match_out565,
   input         match_out566,
   input         match_out567,
   input         match_out568,
   input         match_out569,
   input         match_out570,
   input         match_out571,
   input         match_out572,
   input         match_out573,
   input         match_out574,
   input         match_out575,
   input         match_out576,
   input         match_out577,
   input         match_out578,
   input         match_out579,
   input         match_out580,
   input         match_out581,
   input         match_out582,
   input         match_out583,
   input         match_out584,
   input         match_out585,
   input         match_out586,
   input         match_out587,
   input         match_out588,
   input         match_out589,
   input         match_out590,
   input         match_out591,
   input         match_out592,
   input         match_out593,
   input         match_out594,
   input         match_out595,
   input         match_out596,
   input         match_out597,
   input         match_out598,
   input         match_out599,
   input         match_out600,
   input         match_out601,
   input         match_out602,
   input         match_out603,
   input         match_out604,
   input         match_out605,
   input         match_out606,
   input         match_out607,
   input         match_out608,
   input         match_out609,
   input         match_out610,
   input         match_out611,
   input         match_out612,
   input         match_out613,
   input         match_out614,
   input         match_out615,
   input         match_out616,
   input         match_out617,
   input         match_out618,
   input         match_out619,
   input         match_out620,
   input         match_out621,
   input         match_out622,
   input         match_out623,
   input         match_out624,
   input         match_out625,
   input         match_out626,
   input         match_out627,
   input         match_out628,
   input         match_out629,
   input         match_out630,
   input         match_out631,
   input         match_out632,
   input         match_out633,
   input         match_out634,
   input         match_out635,
   input         match_out636,
   input         match_out637,
   input         match_out638,
   input         match_out639,
   input         match_out640,
   input         match_out641,
   input         match_out642,
   input         match_out643,
   input         match_out644,
   input         match_out645,
   input         match_out646,
   input         match_out647,
   input         match_out648,
   input         match_out649,
   input         match_out650,
   input         match_out651,
   input         match_out652,
   input         match_out653,
   input         match_out654,
   input         match_out655,
   input         match_out656,
   input         match_out657,
   input         match_out658,
   input         match_out659,
   input         match_out660,
   input         match_out661,
   input         match_out662,
   input         match_out663,
   input         match_out664,
   input         match_out665,
   input         match_out666,
   input         match_out667,
   input         match_out668,
   input         match_out669,
   input         match_out670,
   input         match_out671,
   input         match_out672,
   input         match_out673,
   input         match_out674,
   input         match_out675,
   input         match_out676,
   input         match_out677,
   input         match_out678,
   input         match_out679,
   input         match_out680,
   input         match_out681,
   input         match_out682,
   input         match_out683,
   input         match_out684,
   input         match_out685,
   input         match_out686,
   input         match_out687,
   input         match_out688,
   input         match_out689,
   input         match_out690,
   input         match_out691,
   input         match_out692,
   input         match_out693,
   input         match_out694,
   input         match_out695,
   input         match_out696,
   input         match_out697,
   input         match_out698,
   input         match_out699,
   input         match_out700,
   input         match_out701,
   input         match_out702,
   input         match_out703,
   input         match_out704,
   input         match_out705,
   input         match_out706,
   input         match_out707,
   input         match_out708,
   input         match_out709,
   input         match_out710,
   input         match_out711,
   input         match_out712,
   input         match_out713,
   input         match_out714,
   input         match_out715,
   input         match_out716,
   input         match_out717,
   input         match_out718,
   input         match_out719,
   input         match_out720,
   input         match_out721,
   input         match_out722,
   input         match_out723,
   input         match_out724,
   input         match_out725,
   input         match_out726,
   input         match_out727,
   input         match_out728,
   input         match_out729,
   input         match_out730,
   input         match_out731,
   input         match_out732,
   input         match_out733,
   input         match_out734,
   input         match_out735,
   input         match_out736,
   input         match_out737,
   input         match_out738,
   input         match_out739,
   input         match_out740,
   input         match_out741,
   input         match_out742,
   input         match_out743,
   input         match_out744,
   input         match_out745,
   input         match_out746,
   input         match_out747,
   input         match_out748,
   input         match_out749,
   input         match_out750,
   input         match_out751,
   input         match_out752,
   input         match_out753,
   input         match_out754,
   input         match_out755,
   input         match_out756,
   input         match_out757,
   input         match_out758,
   input         match_out759,
   input         match_out760,
   input         match_out761,
   input         match_out762,
   input         match_out763,
   input         match_out764,
   input         match_out765,
   input         match_out766,
   input         match_out767,
   input         match_out768,
   input         match_out769,
   input         match_out770,
   input         match_out771,
   input         match_out772,
   input         match_out773,
   input         match_out774,
   input         match_out775,
   input         match_out776,
   input         match_out777,
   input         match_out778,
   input         match_out779,
   input         match_out780,
   input         match_out781,
   input         match_out782,
   input         match_out783,
   input         match_out784,
   input         match_out785,
   input         match_out786,
   input         match_out787,
   input         match_out788,
   input         match_out789,
   input         match_out790,
   input         match_out791,
   input         match_out792,
   input         match_out793,
   input         match_out794,
   input         match_out795,
   input         match_out796,
   input         match_out797,
   input         match_out798,
   input         match_out799,
   input         match_out800,
   input         match_out801,
   input         match_out802,
   input         match_out803,
   input         match_out804,
   input         match_out805,
   input         match_out806,
   input         match_out807,
   input         match_out808,
   input         match_out809,
   input         match_out810,
   input         match_out811,
   input         match_out812,
   input         match_out813,
   input         match_out814,
   input         match_out815,
   input         match_out816,
   input         match_out817,
   input         match_out818,
   input         match_out819,
   input         match_out820,
   input         match_out821,
   input         match_out822,
   input         match_out823,
   input         match_out824,
   input         match_out825,
   input         match_out826,
   input         match_out827,
   input         match_out828,
   input         match_out829,
   input         match_out830,
   input         match_out831,
   input         match_out832,
   input         match_out833,
   input         match_out834,
   input         match_out835,
   input         match_out836,
   input         match_out837,
   input         match_out838,
   input         match_out839,
   input         match_out840,
   input         match_out841,
   input         match_out842,
   input         match_out843,
   input         match_out844,
   input         match_out845,
   input         match_out846,
   input         match_out847,
   input         match_out848,
   input         match_out849,
   input         match_out850,
   input         match_out851,
   input         match_out852,
   input         match_out853,
   input         match_out854,
   input         match_out855,
   input         match_out856,
   input         match_out857,
   input         match_out858,
   input         match_out859,
   input         match_out860,
   input         match_out861,
   input         match_out862,
   input         match_out863,
   input         match_out864,
   input         match_out865,
   input         match_out866,
   input         match_out867,
   input         match_out868,
   input         match_out869,
   input         match_out870,
   input         match_out871,
   input         match_out872,
   input         match_out873,
   input         match_out874,
   input         match_out875,
   input         match_out876,
   input         match_out877,
   input         match_out878,
   input         match_out879,
   input         match_out880,
   input         match_out881,
   input         match_out882,
   input         match_out883,
   input         match_out884,
   input         match_out885,
   input         match_out886,
   input         match_out887,
   input         match_out888,
   input         match_out889,
   input         match_out890,
   input         match_out891,
   input         match_out892,
   input         match_out893,
   input         match_out894,
   input         match_out895,
   input         match_out896,
   input         match_out897,
   input         match_out898,
   input         match_out899,
   input         match_out900,
   input         match_out901,
   input         match_out902,
   input         match_out903,
   input         match_out904,
   input         match_out905,
   input         match_out906,
   input         match_out907,
   input         match_out908,
   input         match_out909,
   input         match_out910,
   input         match_out911,
   input         match_out912,
   input         match_out913,
   input         match_out914,
   input         match_out915,
   input         match_out916,
   input         match_out917,
   input         match_out918,
   input         match_out919,
   input         match_out920,
   input         match_out921,
   input         match_out922,
   input         match_out923,
   input         match_out924,
   input         match_out925,
   input         match_out926,
   input         match_out927,
   input         match_out928,
   input         match_out929,
   input         match_out930,
   input         match_out931,
   input         match_out932,
   input         match_out933,
   input         match_out934,
   input         match_out935,
   input         match_out936,
   input         match_out937,
   input         match_out938,
   input         match_out939,
   input         match_out940,
   input         match_out941,
   input         match_out942,
   input         match_out943,
   input         match_out944,
   input         match_out945,
   input         match_out946,
   input         match_out947,
   input         match_out948,
   input         match_out949,
   input         match_out950,
   input         match_out951,
   input         match_out952,
   input         match_out953,
   input         match_out954,
   input         match_out955,
   input         match_out956,
   input         match_out957,
   input         match_out958,
   input         match_out959,
   input         match_out960,
   input         match_out961,
   input         match_out962,
   input         match_out963,
   input         match_out964,
   input         match_out965,
   input         match_out966,
   input         match_out967,
   input         match_out968,
   input         match_out969,
   input         match_out970,
   input         match_out971,
   input         match_out972,
   input         match_out973,
   input         match_out974,
   input         match_out975,
   input         match_out976,
   input         match_out977,
   input         match_out978,
   input         match_out979,
   input         match_out980,
   input         match_out981,
   input         match_out982,
   input         match_out983,
   input         match_out984,
   input         match_out985,
   input         match_out986,
   input         match_out987,
   input         match_out988,
   input         match_out989,
   input         match_out990,
   input         match_out991,
   input         match_out992,
   input         match_out993,
   input         match_out994,
   input         match_out995,
   input         match_out996,
   input         match_out997,
   input         match_out998,
   input         match_out999,
   input         match_out1000,
   input         match_out1001,
   input         match_out1002,
   input         match_out1003,
   input         match_out1004,
   input         match_out1005,
   input         match_out1006,
   input         match_out1007,
   input         match_out1008,
   input         match_out1009,
   input         match_out1010,
   input         match_out1011,
   input         match_out1012,
   input         match_out1013,
   input         match_out1014,
   input         match_out1015,
   input         match_out1016,
   input         match_out1017,
   input         match_out1018,
   input         match_out1019,
   input         match_out1020,
   input         match_out1021,
   input         match_out1022,
   input         match_out1023,
   input         match_out1024,
   input         match_out1025,
   input         match_out1026,
   input         match_out1027,
   input         match_out1028,
   input         match_out1029,
   input         match_out1030,
   input         match_out1031,
   input         match_out1032,
   input         match_out1033,
   input         match_out1034,
   input         match_out1035,
   input         match_out1036,
   input         match_out1037,
   input         match_out1038,
   input         match_out1039,
   input         match_out1040,
   input         match_out1041,
   input         match_out1042,
   input         match_out1043,
   input         match_out1044,
   input         match_out1045,
   input         match_out1046,
   input         match_out1047,
   input         match_out1048,
   input         match_out1049,
   input         match_out1050,
   input         match_out1051,
   input         match_out1052,
   input         match_out1053,
   input         match_out1054,
   input         match_out1055,
   input         match_out1056,
   input         match_out1057,
   input         match_out1058,
   input         match_out1059,
   input         match_out1060,
   input         match_out1061,
   input         match_out1062,
   input         match_out1063,
   input         match_out1064,
   input         match_out1065,
   input         match_out1066,
   input         match_out1067,
   input         match_out1068,
   input         match_out1069,
   input         match_out1070,
   input         match_out1071,
   input         match_out1072,
   input         match_out1073,
   input         match_out1074,
   input         match_out1075,
   input         match_out1076,
   input         match_out1077,
   input         match_out1078,
   input         match_out1079,
   input         match_out1080,
   input         match_out1081,
   input         match_out1082,
   input         match_out1083,
   input         match_out1084,
   input         match_out1085,
   input         match_out1086,
   input         match_out1087,
   input         match_out1088,
   input         match_out1089,
   input         match_out1090,
   input         match_out1091,
   input         match_out1092,
   input         match_out1093,
   input         match_out1094,
   input         match_out1095,
   input         match_out1096,
   input         match_out1097,
   input         match_out1098,
   input         match_out1099,
   input         match_out1100,
   input         match_out1101,
   input         match_out1102,
   input         match_out1103,
   input         match_out1104,
   input         match_out1105,
   input         match_out1106,
   input         match_out1107,
   input         match_out1108,
   input         match_out1109,
   input         match_out1110,
   input         match_out1111,
   input         match_out1112,
   input         match_out1113,
   input         match_out1114,
   input         match_out1115,
   input         match_out1116,
   input         match_out1117,
   input         match_out1118,
   input         match_out1119,
   input         match_out1120,
   input         match_out1121,
   input         match_out1122,
   input         match_out1123,
   input         match_out1124,
   input         match_out1125,
   input         match_out1126,
   input         match_out1127,
   input         match_out1128,
   input         match_out1129,
   input         match_out1130,
   input         match_out1131,
   input         match_out1132,
   input         match_out1133,
   input         match_out1134,
   input         match_out1135,
   input         match_out1136,
   input         match_out1137,
   input         match_out1138,
   input         match_out1139,
   input         match_out1140,
   input         match_out1141,
   input         match_out1142,
   input         match_out1143,
   input         match_out1144,
   input         match_out1145,
   input         match_out1146,
   input         match_out1147,
   input         match_out1148,
   input         match_out1149,
   input         match_out1150,
   input         match_out1151,
   input         match_out1152,
   input         match_out1153,
   input         match_out1154,
   input         match_out1155,
   input         match_out1156,
   input         match_out1157,
   input         match_out1158,
   input         match_out1159,
   input         match_out1160,
   input         match_out1161,
   input         match_out1162,
   input         match_out1163,
   input         match_out1164,
   input         match_out1165,
   input         match_out1166,
   input         match_out1167,
   input         match_out1168,
   input         match_out1169,
   input         match_out1170,
   input         match_out1171,
   input         match_out1172,
   input         match_out1173,
   input         match_out1174,
   input         match_out1175,
   input         match_out1176,
   input         match_out1177,
   input         match_out1178,
   input         match_out1179,
   input         match_out1180,
   input         match_out1181,
   input         match_out1182,
   input         match_out1183,
   input         match_out1184,
   input         match_out1185,
   input         match_out1186,
   input         match_out1187,
   input         match_out1188,
   input         match_out1189,
   input         match_out1190,
   input         match_out1191,
   input         match_out1192,
   input         match_out1193,
   input         match_out1194,
   input         match_out1195,
   input         match_out1196,
   input         match_out1197,
   input         match_out1198,
   input         match_out1199,
   input         match_out1200,
   input         match_out1201,
   input         match_out1202,
   input         match_out1203,
   input         match_out1204,
   input         match_out1205,
   input         match_out1206,
   input         match_out1207,
   input         match_out1208,
   input         match_out1209,
   input         match_out1210,
   input         match_out1211,
   input         match_out1212,
   input         match_out1213,
   input         match_out1214,
   input         match_out1215,
   input         match_out1216,
   input         match_out1217,
   input         match_out1218,
   input         match_out1219,
   input         match_out1220,
   input         match_out1221,
   input         match_out1222,
   input         match_out1223,
   input         match_out1224,
   input         match_out1225,
   input         match_out1226,
   input         match_out1227,
   input         match_out1228,
   input         match_out1229,
   input         match_out1230,
   input         match_out1231,
   input         match_out1232,
   input         match_out1233,
   input         match_out1234,
   input         match_out1235,
   input         match_out1236,
   input         match_out1237,
   input         match_out1238,
   input         match_out1239,
   input         match_out1240,
   input         match_out1241,
   input         match_out1242,
   input         match_out1243,
   input         match_out1244,
   input         match_out1245,
   input         match_out1246,
   input         match_out1247,
   input         match_out1248,
   input         match_out1249,
   input         match_out1250,
   input         match_out1251,
   input         match_out1252,
   input         match_out1253,
   input         match_out1254,
   input         match_out1255,
   input         match_out1256,
   input         match_out1257,
   input         match_out1258,
   input         match_out1259,
   input         match_out1260,
   input         match_out1261,
   input         match_out1262,
   input         match_out1263,
   input         match_out1264,
   input         match_out1265,
   input         match_out1266,
   input         match_out1267,
   input         match_out1268,
   input         match_out1269,
   input         match_out1270,
   input         match_out1271,
   input         match_out1272,
   input         match_out1273,
   input         match_out1274,
   input         match_out1275,
   input         match_out1276,
   input         match_out1277,
   input         match_out1278,
   input         match_out1279,
   input         match_out1280,
   input         match_out1281,
   input         match_out1282,
   input         match_out1283,
   input         match_out1284,
   input         match_out1285,
   input         match_out1286,
   input         match_out1287,
   input         match_out1288,
   input         match_out1289,
   input         match_out1290,
   input         match_out1291,
   input         match_out1292,
   input         match_out1293,
   input         match_out1294,
   input         match_out1295,
   input         match_out1296,
   input         match_out1297,
   input         match_out1298,
   input         match_out1299,
   input         match_out1300,
   input         match_out1301,
   input         match_out1302,
   input         match_out1303,
   input         match_out1304,
   input         match_out1305,
   input         match_out1306,
   input         match_out1307,
   input         match_out1308,
   input         match_out1309,
   input         match_out1310,
   input         match_out1311,
   input         match_out1312,
   input         match_out1313,
   input         match_out1314,
   input         match_out1315,
   input         match_out1316,
   input         match_out1317,
   input         match_out1318,
   input         match_out1319,
   input         match_out1320,
   input         match_out1321,
   input         match_out1322,
   input         match_out1323,
   input         match_out1324,
   input         match_out1325,
   input         match_out1326,
   input         match_out1327,
   input         match_out1328,
   input         match_out1329,
   input         match_out1330,
   input         match_out1331,
   input         match_out1332,
   input         match_out1333,
   input         match_out1334,
   input         match_out1335,
   input         match_out1336,
   input         match_out1337,
   input         match_out1338,
   input         match_out1339,
   input         match_out1340,
   input         match_out1341,
   input         match_out1342,
   input         match_out1343,
   input         match_out1344,
   input         match_out1345,
   input         match_out1346,
   input         match_out1347,
   input         match_out1348,
   input         match_out1349,
   input         match_out1350,
   input         match_out1351,
   input         match_out1352,
   input         match_out1353,
   input         match_out1354,
   input         match_out1355,
   input         match_out1356,
   input         match_out1357,
   input         match_out1358,
   input         match_out1359,
   input         match_out1360,
   input         match_out1361,
   input         match_out1362,
   input         match_out1363,
   input         match_out1364,
   input         match_out1365,
   input         match_out1366,
   input         match_out1367,
   input         match_out1368,
   input         match_out1369,
   input         match_out1370,
   input         match_out1371,
   input         match_out1372,
   input         match_out1373,
   input         match_out1374,
   input         match_out1375,
   input         match_out1376,
   input         match_out1377,
   input         match_out1378,
   input         match_out1379,
   input         match_out1380,
   input         match_out1381,
   input         match_out1382,
   input         match_out1383,
   input         match_out1384,
   input         match_out1385,
   input         match_out1386,
   input         match_out1387,
   input         match_out1388,
   input         match_out1389,
   input         match_out1390,
   input         match_out1391,
   input         match_out1392,
   input         match_out1393,
   input         match_out1394,
   input         match_out1395,
   input         match_out1396,
   input         match_out1397,
   input         match_out1398,
   input         match_out1399,
   input         match_out1400,
   input         match_out1401,
   input         match_out1402,
   input         match_out1403,
   input         match_out1404,
   input         match_out1405,
   input         match_out1406,
   input         match_out1407,
   input         match_out1408,
   input         match_out1409,
   input         match_out1410,
   input         match_out1411,
   input         match_out1412,
   input         match_out1413,
   input         match_out1414,
   input         match_out1415,
   input         match_out1416,
   input         match_out1417,
   input         match_out1418,
   input         match_out1419,
   input         match_out1420,
   input         match_out1421,
   input         match_out1422,
   input         match_out1423,
   input         match_out1424,
   input         match_out1425,
   input         match_out1426,
   input         match_out1427,
   input         match_out1428,
   input         match_out1429,
   input         match_out1430,
   input         match_out1431,
   input         match_out1432,
   input         match_out1433,
   input         match_out1434,
   input         match_out1435,
   input         match_out1436,
   input         match_out1437,
   input         match_out1438,
   input         match_out1439,
   input         match_out1440,
   input         match_out1441,
   input         match_out1442,
   input         match_out1443,
   input         match_out1444,
   input         match_out1445,
   input         match_out1446,
   input         match_out1447,
   input         match_out1448,
   input         match_out1449,
   input         match_out1450,
   input         match_out1451,
   input         match_out1452,
   input         match_out1453,
   input         match_out1454,
   input         match_out1455,
   input         match_out1456,
   input         match_out1457,
   input         match_out1458,
   input         match_out1459,
   input         match_out1460,
   input         match_out1461,
   input         match_out1462,
   input         match_out1463,
   input         match_out1464,
   input         match_out1465,
   input         match_out1466,
   input         match_out1467,
   input         match_out1468,
   input         match_out1469,
   input         match_out1470,
   input         match_out1471,
   input         match_out1472,
   input         match_out1473,
   input         match_out1474,
   input         match_out1475,
   input         match_out1476,
   input         match_out1477,
   input         match_out1478,
   input         match_out1479,
   input         match_out1480,
   input         match_out1481,
   input         match_out1482,
   input         match_out1483,
   input         match_out1484,
   input         match_out1485,
   input         match_out1486,
   input         match_out1487,
   input         match_out1488,
   input         match_out1489,
   input         match_out1490,
   input         match_out1491,
   input         match_out1492,
   input         match_out1493,
   input         match_out1494,
   input         match_out1495,
   input         match_out1496,
   input         match_out1497,
   input         match_out1498,
   input         match_out1499,
   input         match_out1500,
   input         match_out1501,
   input         match_out1502,
   input         match_out1503,
   input         match_out1504,
   input         match_out1505,
   input         match_out1506,
   input         match_out1507,
   input         match_out1508,
   input         match_out1509,
   input         match_out1510,
   input         match_out1511,
   input         match_out1512,
   input         match_out1513,
   input         match_out1514,
   input         match_out1515,
   input         match_out1516,
   input         match_out1517,
   input         match_out1518,
   input         match_out1519,
   input         match_out1520,
   input         match_out1521,
   input         match_out1522,
   input         match_out1523,
   input         match_out1524,
   input         match_out1525,
   input         match_out1526,
   input         match_out1527,
   input         match_out1528,
   input         match_out1529,
   input         match_out1530,
   input         match_out1531,
   input         match_out1532,
   input         match_out1533,
   input         match_out1534,
   input         match_out1535,
   input         match_out1536,
   input         match_out1537,
   input         match_out1538,
   input         match_out1539,
   input         match_out1540,
   input         match_out1541,
   input         match_out1542,
   input         match_out1543,
   input         match_out1544,
   input         match_out1545,
   input         match_out1546,
   input         match_out1547,
   input         match_out1548,
   input         match_out1549,
   input         match_out1550,
   input         match_out1551,
   input         match_out1552,
   input         match_out1553,
   input         match_out1554,
   input         match_out1555,
   input         match_out1556,
   input         match_out1557,
   input         match_out1558,
   input         match_out1559,
   input         match_out1560,
   input         match_out1561,
   input         match_out1562,
   input         match_out1563,
   input         match_out1564,
   input         match_out1565,
   input         match_out1566,
   input         match_out1567,
   input         match_out1568,
   input         match_out1569,
   input         match_out1570,
   input         match_out1571,
   input         match_out1572,
   input         match_out1573,
   input         match_out1574,
   input         match_out1575,
   input         match_out1576,
   input         match_out1577,
   input         match_out1578,
   input         match_out1579,
   input         match_out1580,
   input         match_out1581,
   input         match_out1582,
   input         match_out1583,
   input         match_out1584,
   input         match_out1585,
   input         match_out1586,
   input         match_out1587,
   input         match_out1588,
   input         match_out1589,
   input         match_out1590,
   input         match_out1591,
   input         match_out1592,
   input         match_out1593,
   input         match_out1594,
   input         match_out1595,
   input         match_out1596,
   input         match_out1597,
   input         match_out1598,
   input         match_out1599,
   input         match_out1600,
   input         match_out1601,
   input         match_out1602,
   input         match_out1603,
   input         match_out1604,
   input         match_out1605,
   input         match_out1606,
   input         match_out1607,
   input         match_out1608,
   input         match_out1609,
   input         match_out1610,
   input         match_out1611,
   input         match_out1612,
   input         match_out1613,
   input         match_out1614,
   input         match_out1615,
   input         match_out1616,
   input         match_out1617,
   input         match_out1618,
   input         match_out1619,
   input         match_out1620,
   input         match_out1621,
   input         match_out1622,
   input         match_out1623,
   input         match_out1624,
   input         match_out1625,
   input         match_out1626,
   input         match_out1627,
   input         match_out1628,
   input         match_out1629,
   input         match_out1630,
   input         match_out1631,
   input         match_out1632,
   input         match_out1633,
   input         match_out1634,
   input         match_out1635,
   input         match_out1636,
   input         match_out1637,
   input         match_out1638,
   input         match_out1639,
   input         match_out1640,
   input         match_out1641,
   input         match_out1642,
   input         match_out1643,
   input         match_out1644,
   input         match_out1645,
   input         match_out1646,
   input         match_out1647,
   input         match_out1648,
   input         match_out1649,
   input         match_out1650,
   input         match_out1651,
   input         match_out1652,
   input         match_out1653,
   input         match_out1654,
   input         match_out1655,
   input         match_out1656,
   input         match_out1657,
   input         match_out1658,
   input         match_out1659,
   input         match_out1660,
   input         match_out1661,
   input         match_out1662,
   input         match_out1663,
   input         match_out1664,
   input         match_out1665,
   input         match_out1666,
   input         match_out1667,
   input         match_out1668,
   input         match_out1669,
   input         match_out1670,
   input         match_out1671,
   input         match_out1672,
   input         match_out1673,
   input         match_out1674,
   input         match_out1675,
   input         match_out1676,
   input         match_out1677,
   input         match_out1678,
   input         match_out1679,
   input         match_out1680,
   input         match_out1681,
   input         match_out1682,
   input         match_out1683,
   input         match_out1684,
   input         match_out1685,
   input         match_out1686,
   input         match_out1687,
   input         match_out1688,
   input         match_out1689,
   input         match_out1690,
   input         match_out1691,
   input         match_out1692,
   input         match_out1693,
   input         match_out1694,
   input         match_out1695,
   input         match_out1696,
   input         match_out1697,
   input         match_out1698,
   input         match_out1699,
   input         match_out1700,
   input         match_out1701,
   input         match_out1702,
   input         match_out1703,
   input         match_out1704,
   input         match_out1705,
   input         match_out1706,
   input         match_out1707,
   input         match_out1708,
   input         match_out1709,
   input         match_out1710,
   input         match_out1711,
   input         match_out1712,
   input         match_out1713,
   input         match_out1714,
   input         match_out1715,
   input         match_out1716,
   input         match_out1717,
   input         match_out1718,
   input         match_out1719,
   input         match_out1720,
   input         match_out1721,
   input         match_out1722,
   input         match_out1723,
   input         match_out1724,
   input         match_out1725,
   input         match_out1726,
   input         match_out1727,
   input         match_out1728,
   input         match_out1729,
   input         match_out1730,
   input         match_out1731,
   input         match_out1732,
   input         match_out1733,
   input         match_out1734,
   input         match_out1735,
   input         match_out1736,
   input         match_out1737,
   input         match_out1738,
   input         match_out1739,
   input         match_out1740,
   input         match_out1741,
   input         match_out1742,
   input         match_out1743,
   input         match_out1744,
   input         match_out1745,
   input         match_out1746,
   input         match_out1747,
   input         match_out1748,
   input         match_out1749,
   input         match_out1750,
   input         match_out1751,
   input         match_out1752,
   input         match_out1753,
   input         match_out1754,
   input         match_out1755,
   input         match_out1756,
   input         match_out1757,
   input         match_out1758,
   input         match_out1759,
   input         match_out1760,
   input         match_out1761,
   input         match_out1762,
   input         match_out1763,
   input         match_out1764,
   input         match_out1765,
   input         match_out1766,
   input         match_out1767,
   input         match_out1768,
   input         match_out1769,
   input         match_out1770,
   input         match_out1771,
   input         match_out1772,
   input         match_out1773,
   input         match_out1774,
   input         match_out1775,
   input         match_out1776,
   input         match_out1777,
   input         match_out1778,
   input         match_out1779,
   input         match_out1780,
   input         match_out1781,
   input         match_out1782,
   input         match_out1783,
   input         match_out1784,
   input         match_out1785,
   input         match_out1786,
   input         match_out1787,
   input         match_out1788,
   input         match_out1789,
   input         match_out1790,
   input         match_out1791,
   input         match_out1792,
   input         match_out1793,
   input         match_out1794,
   input         match_out1795,
   input         match_out1796,
   input         match_out1797,
   input         match_out1798,
   input         match_out1799,
   input         match_out1800,
   input         match_out1801,
   input         match_out1802,
   input         match_out1803,
   input         match_out1804,
   input         match_out1805,
   input         match_out1806,
   input         match_out1807,
   input         match_out1808,
   input         match_out1809,
   input         match_out1810,
   input         match_out1811,
   input         match_out1812,
   input         match_out1813,
   input         match_out1814,
   input         match_out1815,
   input         match_out1816,
   input         match_out1817,
   input         match_out1818,
   input         match_out1819,
   input         match_out1820,
   input         match_out1821,
   input         match_out1822,
   input         match_out1823,
   input         match_out1824,
   input         match_out1825,
   input         match_out1826,
   input         match_out1827,
   input         match_out1828,
   input         match_out1829,
   input         match_out1830,
   input         match_out1831,
   input         match_out1832,
   input         match_out1833,
   input         match_out1834,
   input         match_out1835,
   input         match_out1836,
   input         match_out1837,
   input         match_out1838,
   input         match_out1839,
   input         match_out1840,
   input         match_out1841,
   input         match_out1842,
   input         match_out1843,
   input         match_out1844,
   input         match_out1845,
   input         match_out1846,
   input         match_out1847,
   input         match_out1848,
   input         match_out1849,
   input         match_out1850,
   input         match_out1851,
   input         match_out1852,
   input         match_out1853,
   input         match_out1854,
   input         match_out1855,
   input         match_out1856,
   input         match_out1857,
   input         match_out1858,
   input         match_out1859,
   input         match_out1860,
   input         match_out1861,
   input         match_out1862,
   input         match_out1863,
   input         match_out1864,
   input         match_out1865,
   input         match_out1866,
   input         match_out1867,
   input         match_out1868,
   input         match_out1869,
   input         match_out1870,
   input         match_out1871,
   input         match_out1872,
   input         match_out1873,
   input         match_out1874,
   input         match_out1875,
   input         match_out1876,
   input         match_out1877,
   input         match_out1878,
   input         match_out1879,
   input         match_out1880,
   input         match_out1881,
   input         match_out1882,
   input         match_out1883,
   input         match_out1884,
   input         match_out1885,
   input         match_out1886,
   input         match_out1887,
   input         match_out1888,
   input         match_out1889,
   input         match_out1890,
   input         match_out1891,
   input         match_out1892,
   input         match_out1893,
   input         match_out1894,
   input         match_out1895,
   input         match_out1896,
   input         match_out1897,
   input         match_out1898,
   input         match_out1899,
   input         match_out1900,
   input         match_out1901,
   input         match_out1902,
   input         match_out1903,
   input         match_out1904,
   input         match_out1905,
   input         match_out1906,
   input         match_out1907,
   input         match_out1908,
   input         match_out1909,
   input         match_out1910,
   input         match_out1911,
   input         match_out1912,
   input         match_out1913,
   input         match_out1914,
   input         match_out1915,
   input         match_out1916,
   input         match_out1917,
   input         match_out1918,
   input         match_out1919,
   input         match_out1920,
   input         match_out1921,
   input         match_out1922,
   input         match_out1923,
   input         match_out1924,
   input         match_out1925,
   input         match_out1926,
   input         match_out1927,
   input         match_out1928,
   input         match_out1929,
   input         match_out1930,
   input         match_out1931,
   input         match_out1932,
   input         match_out1933,
   input         match_out1934,
   input         match_out1935,
   input         match_out1936,
   input         match_out1937,
   input         match_out1938,
   input         match_out1939,
   input         match_out1940,
   input         match_out1941,
   input         match_out1942,
   input         match_out1943,
   input         match_out1944,
   input         match_out1945,
   input         match_out1946,
   input         match_out1947,
   input         match_out1948,
   input         match_out1949,
   input         match_out1950,
   input         match_out1951,
   input         match_out1952,
   input         match_out1953,
   input         match_out1954,
   input         match_out1955,
   input         match_out1956,
   input         match_out1957,
   input         match_out1958,
   input         match_out1959,
   input         match_out1960,
   input         match_out1961,
   input         match_out1962,
   input         match_out1963,
   input         match_out1964,
   input         match_out1965,
   input         match_out1966,
   input         match_out1967,
   input         match_out1968,
   input         match_out1969,
   input         match_out1970,
   input         match_out1971,
   input         match_out1972,
   input         match_out1973,
   input         match_out1974,
   input         match_out1975,
   input         match_out1976,
   input         match_out1977,
   input         match_out1978,
   input         match_out1979,
   input         match_out1980,
   input         match_out1981,
   input         match_out1982,
   input         match_out1983,
   input         match_out1984,
   input         match_out1985,
   input         match_out1986,
   input         match_out1987,
   input         match_out1988,
   input         match_out1989,
   input         match_out1990,
   input         match_out1991,
   input         match_out1992,
   input         match_out1993,
   input         match_out1994,
   input         match_out1995,
   input         match_out1996,
   input         match_out1997,
   input         match_out1998,
   input         match_out1999,
   input         match_out2000,
   input         match_out2001,
   input         match_out2002,
   input         match_out2003,
   input         match_out2004,
   input         match_out2005,
   input         match_out2006,
   input         match_out2007,
   input         match_out2008,
   input         match_out2009,
   input         match_out2010,
   input         match_out2011,
   input         match_out2012,
   input         match_out2013,
   input         match_out2014,
   input         match_out2015,
   input         match_out2016,
   input         match_out2017,
   input         match_out2018,
   input         match_out2019,
   input         match_out2020,
   input         match_out2021,
   input         match_out2022,
   input         match_out2023,
   input         match_out2024,
   input         match_out2025,
   input         match_out2026,
   input         match_out2027,
   input         match_out2028,
   input         match_out2029,
   input         match_out2030,
   input         match_out2031,
   input         match_out2032,
   input         match_out2033,
   input         match_out2034,
   input         match_out2035,
   input         match_out2036,
   input         match_out2037,
   input         match_out2038,
   input         match_out2039,
   input         match_out2040,
   input         match_out2041,
   input         match_out2042,
   input         match_out2043,
   input         match_out2044,
   input         match_out2045,
   input         match_out2046,
   input         match_out2047,
   input         match_out2048,
   input         match_out2049,
   input         match_out2050,
   input         match_out2051,
   input         match_out2052,
   input         match_out2053,
   input         match_out2054,
   input         match_out2055,
   input         match_out2056,
   input         match_out2057,
   input         match_out2058,
   input         match_out2059,
   input         match_out2060,
   input         match_out2061,
   input         match_out2062,
   input         match_out2063,
   input         match_out2064,
   input         match_out2065,
   input         match_out2066,
   input         match_out2067,
   input         match_out2068,
   input         match_out2069,
   input         match_out2070,
   input         match_out2071,
   input         match_out2072,
   input         match_out2073,
   input         match_out2074,
   input         match_out2075,
   input         match_out2076,
   input         match_out2077,
   input         match_out2078,
   input         match_out2079,
   input         match_out2080,
   input         match_out2081,
   input         match_out2082,
   input         match_out2083,
   input         match_out2084,
   input         match_out2085,
   input         match_out2086,
   input         match_out2087,
   input         match_out2088,
   input         match_out2089,
   input         match_out2090,
   input         match_out2091,
   input         match_out2092,
   input         match_out2093,
   input         match_out2094,
   input         match_out2095,
   input         match_out2096,
   input         match_out2097,
   input         match_out2098,
   input         match_out2099,
   input         match_out2100,
   input         match_out2101,
   input         match_out2102,
   input         match_out2103,
   input         match_out2104,
   input         match_out2105,
   input         match_out2106,
   input         match_out2107,
   input         match_out2108,
   input         match_out2109,
   input         match_out2110,
   input         match_out2111,
   input         match_out2112,
   input         match_out2113,
   input         match_out2114,
   input         match_out2115,
   input         match_out2116,
   input         match_out2117,
   input         match_out2118,
   input         match_out2119,
   input         match_out2120,
   input         match_out2121,
   input         match_out2122,
   input         match_out2123,
   input         match_out2124,
   input         match_out2125,
   input         match_out2126,
   input         match_out2127,
   input         match_out2128,
   input         match_out2129,
   input         match_out2130,
   input         match_out2131,
   input         match_out2132,
   input         match_out2133,
   input         match_out2134,
   input         match_out2135,
   input         match_out2136,
   input         match_out2137,
   input         match_out2138,
   input         match_out2139,
   input         match_out2140,
   input         match_out2141,
   input         match_out2142,
   input         match_out2143,
   input         match_out2144,
   input         match_out2145,
   input         match_out2146,
   input         match_out2147,
   input         match_out2148,
   input         match_out2149,
   input         match_out2150,
   input         match_out2151,
   input         match_out2152,
   input         match_out2153,
   input         match_out2154,
   input         match_out2155,
   input         match_out2156,
   input         match_out2157,
   input         match_out2158,
   input         match_out2159,
   input         match_out2160,
   input         match_out2161,
   input         match_out2162,
   input         match_out2163,
   input         match_out2164,
   input         match_out2165,
   input         match_out2166,
   input         match_out2167,
   input         match_out2168,
   input         match_out2169,
   input         match_out2170,
   input         match_out2171,
   input         match_out2172,
   input         match_out2173,
   input         match_out2174,
   input         match_out2175,
   input         match_out2176,
   input         match_out2177,
   input         match_out2178,
   input         match_out2179,
   input         match_out2180,
   input         match_out2181,
   input         match_out2182,
   input         match_out2183,
   input         match_out2184,
   input         match_out2185,
   input         match_out2186,
   input         match_out2187,
   input         match_out2188,
   input         match_out2189,
   input         match_out2190,
   input         match_out2191,
   input         match_out2192,
   input         match_out2193,
   input         match_out2194,
   input         match_out2195,
   input         match_out2196,
   input         match_out2197,
   input         match_out2198,
   input         match_out2199,
   input         match_out2200,
   input         match_out2201,
   input         match_out2202,
   input         match_out2203,
   input         match_out2204,
   input         match_out2205,
   input         match_out2206,
   input         match_out2207,
   input         match_out2208,
   input         match_out2209,
   input         match_out2210,
   input         match_out2211,
   input         match_out2212,
   input         match_out2213,
   input         match_out2214,
   input         match_out2215,
   input         match_out2216,
   input         match_out2217,
   input         match_out2218,
   input         match_out2219,
   input         match_out2220,
   input         match_out2221,
   input         match_out2222,
   input         match_out2223,
   input         match_out2224,
   input         match_out2225,
   input         match_out2226,
   input         match_out2227,
   input         match_out2228,
   input         match_out2229,
   input         match_out2230,
   input         match_out2231,
   input         match_out2232,
   input         match_out2233,
   input         match_out2234,
   input         match_out2235,
   input         match_out2236,
   input         match_out2237,
   input         match_out2238,
   input         match_out2239,
   input         match_out2240,
   input         match_out2241,
   input         match_out2242,
   input         match_out2243,
   input         match_out2244,
   input         match_out2245,
   input         match_out2246,
   input         match_out2247,
   input         match_out2248,
   input         match_out2249,
   input         match_out2250,
   input         match_out2251,
   input         match_out2252,
   input         match_out2253,
   input         match_out2254,
   input         match_out2255,
   input         match_out2256,
   input         match_out2257,
   input         match_out2258,
   input         match_out2259,
   input         match_out2260,
   input         match_out2261,
   input         match_out2262,
   input         match_out2263,
   input         match_out2264,
   input         match_out2265,
   input         match_out2266,
   input         match_out2267,
   input         match_out2268,
   input         match_out2269,
   input         match_out2270,
   input         match_out2271,
   input         match_out2272,
   input         match_out2273,
   input         match_out2274,
   input         match_out2275,
   input         match_out2276,
   input         match_out2277,
   input         match_out2278,
   input         match_out2279,
   input         match_out2280,
   input         match_out2281,
   input         match_out2282,
   input         match_out2283,
   input         match_out2284,
   input         match_out2285,
   input         match_out2286,
   input         match_out2287,
   input         match_out2288,
   input         match_out2289,
   input         match_out2290,
   input         match_out2291,
   input         match_out2292,
   input         match_out2293,
   input         match_out2294,
   input         match_out2295,
   input         match_out2296,
   input         match_out2297,
   input         match_out2298,
   input         match_out2299,
   input         match_out2300,
   input         match_out2301,
   input         match_out2302,
   input         match_out2303,
   input         match_out2304,
   input         match_out2305,
   input         match_out2306,
   input         match_out2307,
   input         match_out2308,
   input         match_out2309,
   input         match_out2310,
   input         match_out2311,
   input         match_out2312,
   input         match_out2313,
   input         match_out2314,
   input         match_out2315,
   input         match_out2316,
   input         match_out2317,
   input         match_out2318,
   input         match_out2319,
   input         match_out2320,
   input         match_out2321,
   input         match_out2322,
   input         match_out2323,
   input         match_out2324,
   input         match_out2325,
   input         match_out2326,
   input         match_out2327,
   input         match_out2328,
   input         match_out2329,
   input         match_out2330,
   input         match_out2331,
   input         match_out2332,
   input         match_out2333,
   input         match_out2334,
   input         match_out2335,
   input         match_out2336,
   input         match_out2337,
   input         match_out2338,
   input         match_out2339,
   input         match_out2340,
   input         match_out2341,
   input         match_out2342,
   input         match_out2343,
   input         match_out2344,
   input         match_out2345,
   input         match_out2346,
   input         match_out2347,
   input         match_out2348,
   input         match_out2349,
   input         match_out2350,
   input         match_out2351,
   input         match_out2352,
   input         match_out2353,
   input         match_out2354,
   input         match_out2355,
   input         match_out2356,
   input         match_out2357,
   input         match_out2358,
   input         match_out2359,
   input         match_out2360,
   input         match_out2361,
   input         match_out2362,
   input         match_out2363,
   input         match_out2364,
   input         match_out2365,
   input         match_out2366,
   input         match_out2367,
   input         match_out2368,
   input         match_out2369,
   input         match_out2370,
   input         match_out2371,
   input         match_out2372,
   input         match_out2373,
   input         match_out2374,
   input         match_out2375,
   input         match_out2376,
   input         match_out2377,
   input         match_out2378,
   input         match_out2379,
   input         match_out2380,
   input         match_out2381,
   input         match_out2382,
   input         match_out2383,
   input         match_out2384,
   input         match_out2385,
   input         match_out2386,
   input         match_out2387,
   input         match_out2388,
   input         match_out2389,
   input         match_out2390,
   input         match_out2391,
   input         match_out2392,
   input         match_out2393,
   input         match_out2394,
   input         match_out2395,
   input         match_out2396,
   input         match_out2397,
   input         match_out2398,
   input         match_out2399,
   input         match_out2400,
   input         match_out2401,
   input         match_out2402,
   input         match_out2403,
   input         match_out2404,
   input         match_out2405,
   input         match_out2406,
   input         match_out2407,
   input         match_out2408,
   input         match_out2409,
   input         match_out2410,
   input         match_out2411,
   input         match_out2412,
   input         match_out2413,
   input         match_out2414,
   input         match_out2415,
   input         match_out2416,
   input         match_out2417,
   input         match_out2418,
   input         match_out2419,
   input         match_out2420,
   input         match_out2421,
   input         match_out2422,
   input         match_out2423,
   input         match_out2424,
   input         match_out2425,
   input         match_out2426,
   input         match_out2427,
   input         match_out2428,
   input         match_out2429,
   input         match_out2430,
   input         match_out2431,
   input         match_out2432,
   input         match_out2433,
   input         match_out2434,
   input         match_out2435,
   input         match_out2436,
   input         match_out2437,
   input         match_out2438,
   input         match_out2439,
   input         match_out2440,
   input         match_out2441,
   input         match_out2442,
   input         match_out2443,
   input         match_out2444,
   input         match_out2445,
   input         match_out2446,
   input         match_out2447,
   input         match_out2448,
   input         match_out2449,
   input         match_out2450,
   input         match_out2451,
   input         match_out2452,
   input         match_out2453,
   input         match_out2454,
   input         match_out2455,
   input         match_out2456,
   input         match_out2457,
   input         match_out2458,
   input         match_out2459,
   input         match_out2460,
   input         match_out2461,
   input         match_out2462,
   input         match_out2463,
   input         match_out2464,
   input         match_out2465,
   input         match_out2466,
   input         match_out2467,
   input         match_out2468,
   input         match_out2469,
   input         match_out2470,
   input         match_out2471,
   input         match_out2472,
   input         match_out2473,
   input         match_out2474,
   input         match_out2475,
   input         match_out2476,
   input         match_out2477,
   input         match_out2478,
   input         match_out2479,
   input         match_out2480,
   input         match_out2481,
   input         match_out2482,
   input         match_out2483,
   input         match_out2484,
   input         match_out2485,
   input         match_out2486,
   input         match_out2487,
   input         match_out2488,
   input         match_out2489,
   input         match_out2490,
   input         match_out2491,
   input         match_out2492,
   input         match_out2493,
   input         match_out2494,
   input         match_out2495,
   input         match_out2496,
   input         match_out2497,
   input         match_out2498,
   input         match_out2499,
   input         match_out2500,
   input         match_out2501,
   input         match_out2502,
   input         match_out2503,
   input         match_out2504,
   input         match_out2505,
   input         match_out2506,
   input         match_out2507,
   input         match_out2508,
   input         match_out2509,
   input         match_out2510,
   input         match_out2511,
   input         match_out2512,
   input         match_out2513,
   input         match_out2514,
   input         match_out2515,
   input         match_out2516,
   input         match_out2517,
   input         match_out2518,
   input         match_out2519,
   input         match_out2520,
   input         match_out2521,
   input         match_out2522,
   input         match_out2523,
   input         match_out2524,
   input         match_out2525,
   input         match_out2526,
   input         match_out2527,
   input         match_out2528,
   input         match_out2529,
   input         match_out2530,
   input         match_out2531,
   input         match_out2532,
   input         match_out2533,
   input         match_out2534,
   input         match_out2535,
   input         match_out2536,
   input         match_out2537,
   input         match_out2538,
   input         match_out2539,
   input         match_out2540,
   input         match_out2541,
   input         match_out2542,
   input         match_out2543,
   input         match_out2544,
   input         match_out2545,
   input         match_out2546,
   input         match_out2547,
   input         match_out2548,
   input         match_out2549,
   input         match_out2550,
   input         match_out2551,
   input         match_out2552,
   input         match_out2553,
   input         match_out2554,
   input         match_out2555,
   input         match_out2556,
   input         match_out2557,
   input         match_out2558,
   input         match_out2559,
   input         match_out2560,
   input         match_out2561,
   input         match_out2562,
   input         match_out2563,
   input         match_out2564,
   input         match_out2565,
   input         match_out2566,
   input         match_out2567,
   input         match_out2568,
   input         match_out2569,
   input         match_out2570,
   input         match_out2571,
   input         match_out2572,
   input         match_out2573,
   input         match_out2574,
   input         match_out2575,
   input         match_out2576,
   input         match_out2577,
   input         match_out2578,
   input         match_out2579,
   input         match_out2580,
   input         match_out2581,
   input         match_out2582,
   input         match_out2583,
   input         match_out2584,
   input         match_out2585,
   input         match_out2586,
   input         match_out2587,
   input         match_out2588,
   input         match_out2589,
   input         match_out2590,
   input         match_out2591,
   input         match_out2592,
   input         match_out2593,
   input         match_out2594,
   input         match_out2595,
   input         match_out2596,
   input         match_out2597,
   input         match_out2598,
   input         match_out2599,
   input         match_out2600,
   input         match_out2601,
   input         match_out2602,
   input         match_out2603,
   input         match_out2604,
   input         match_out2605,
   input         match_out2606,
   input         match_out2607,
   input         match_out2608,
   input         match_out2609,
   input         match_out2610,
   input         match_out2611,
   input         match_out2612,
   input         match_out2613,
   input         match_out2614,
   input         match_out2615,
   input         match_out2616,
   input         match_out2617,
   input         match_out2618,
   input         match_out2619,
   input         match_out2620,
   input         match_out2621,
   input         match_out2622,
   input         match_out2623,
   input         match_out2624,
   input         match_out2625,
   input         match_out2626,
   input         match_out2627,
   input         match_out2628,
   input         match_out2629,
   input         match_out2630,
   input         match_out2631,
   input         match_out2632,
   input         match_out2633,
   input         match_out2634,
   input         match_out2635,
   input         match_out2636,
   input         match_out2637,
   input         match_out2638,
   input         match_out2639,
   input         match_out2640,
   input         match_out2641,
   input         match_out2642,
   input         match_out2643,
   input         match_out2644,
   input         match_out2645,
   input         match_out2646,
   input         match_out2647,
   input         match_out2648,
   input         match_out2649,
   input         match_out2650,
   input         match_out2651,
   input         match_out2652,
   input         match_out2653,
   input         match_out2654,
   input         match_out2655,
   input         match_out2656,
   input         match_out2657,
   input         match_out2658,
   input         match_out2659,
   input         match_out2660,
   input         match_out2661,
   input         match_out2662,
   input         match_out2663,
   input         match_out2664,
   input         match_out2665,
   input         match_out2666,
   input         match_out2667,
   input         match_out2668,
   input         match_out2669,
   input         match_out2670,
   input         match_out2671,
   input         match_out2672,
   input         match_out2673,
   input         match_out2674,
   input         match_out2675,
   input         match_out2676,
   input         match_out2677,
   input         match_out2678,
   input         match_out2679,
   input         match_out2680,
   input         match_out2681,
   input         match_out2682,
   input         match_out2683,
   input         match_out2684,
   input         match_out2685,
   input         match_out2686,
   input         match_out2687,
   input         match_out2688,
   input         match_out2689,
   input         match_out2690,
   input         match_out2691,
   input         match_out2692,
   input         match_out2693,
   input         match_out2694,
   input         match_out2695,
   input         match_out2696,
   input         match_out2697,
   input         match_out2698,
   input         match_out2699,
   input         match_out2700,
   input         match_out2701,
   input         match_out2702,
   input         match_out2703,
   input         match_out2704,
   input         match_out2705,
   input         match_out2706,
   input         match_out2707,
   input         match_out2708,
   input         match_out2709,
   input         match_out2710,
   input         match_out2711,
   input         match_out2712,
   input         match_out2713,
   input         match_out2714,
   input         match_out2715,
   input         match_out2716,
   input         match_out2717,
   input         match_out2718,
   input         match_out2719,
   input         match_out2720,
   input         match_out2721,
   input         match_out2722,
   input         match_out2723,
   input         match_out2724,
   input         match_out2725,
   input         match_out2726,
   input         match_out2727,
   input         match_out2728,
   input         match_out2729,
   input         match_out2730,
   input         match_out2731,
   input         match_out2732,
   input         match_out2733,
   input         match_out2734,
   input         match_out2735,
   input         match_out2736,
   input         match_out2737,
   input         match_out2738,
   input         match_out2739,
   input         match_out2740,
   input         match_out2741,
   input         match_out2742,
   input         match_out2743,
   input         match_out2744,
   input         match_out2745,
   input         match_out2746,
   input         match_out2747,
   input         match_out2748,
   input         match_out2749,
   input         match_out2750,
   input         match_out2751,
   input         match_out2752,
   input         match_out2753,
   input         match_out2754,
   input         match_out2755,
   input         match_out2756,
   input         match_out2757,
   input         match_out2758,
   input         match_out2759,
   input         match_out2760,
   input         match_out2761,
   input         match_out2762,
   input         match_out2763,
   input         match_out2764,
   input         match_out2765,
   input         match_out2766,
   input         match_out2767,
   input         match_out2768,
   input         match_out2769,
   input         match_out2770,
   input         match_out2771,
   input         match_out2772,
   input         match_out2773,
   input         match_out2774,
   input         match_out2775,
   input         match_out2776,
   input         match_out2777,
   input         match_out2778,
   input         match_out2779,
   input         match_out2780,
   input         match_out2781,
   input         match_out2782,
   input         match_out2783,
   input         match_out2784,
   input         match_out2785,
   input         match_out2786,
   input         match_out2787,
   input         match_out2788,
   input         match_out2789,
   input         match_out2790,
   input         match_out2791,
   input         match_out2792,
   input         match_out2793,
   input         match_out2794,
   input         match_out2795,
   input         match_out2796,
   input         match_out2797,
   input         match_out2798,
   input         match_out2799,
   input         match_out2800,
   input         match_out2801,
   input         match_out2802,
   input         match_out2803,
   input         match_out2804,
   input         match_out2805,
   input         match_out2806,
   input         match_out2807,
   input         match_out2808,
   input         match_out2809,
   input         match_out2810,
   input         match_out2811,
   input         match_out2812,
   input         match_out2813,
   input         match_out2814,
   input         match_out2815,
   input         match_out2816,
   input         match_out2817,
   input         match_out2818,
   input         match_out2819,
   input         match_out2820,
   input         match_out2821,
   input         match_out2822,
   input         match_out2823,
   input         match_out2824,
   input         match_out2825,
   input         match_out2826,
   input         match_out2827,
   input         match_out2828,
   input         match_out2829,
   input         match_out2830,
   input         match_out2831,
   input         match_out2832,
   input         match_out2833,
   input         match_out2834,
   input         match_out2835,
   input         match_out2836,
   input         match_out2837,
   input         match_out2838,
   input         match_out2839,
   input         match_out2840,
   input         match_out2841,
   input         match_out2842,
   input         match_out2843,
   input         match_out2844,
   input         match_out2845,
   input         match_out2846,
   input         match_out2847,
   input         match_out2848,
   input         match_out2849,
   input         match_out2850,
   input         match_out2851,
   input         match_out2852,
   input         match_out2853,
   input         match_out2854,
   input         match_out2855,
   input         match_out2856,
   input         match_out2857,
   input         match_out2858,
   input         match_out2859,
   input         match_out2860,
   input         match_out2861,
   input         match_out2862,
   input         match_out2863,
   input         match_out2864,
   input         match_out2865,
   input         match_out2866,
   input         match_out2867,
   input         match_out2868,
   input         match_out2869,
   input         match_out2870,
   input         match_out2871,
   input         match_out2872,
   input         match_out2873,
   input         match_out2874,
   input         match_out2875,
   input         match_out2876,
   input         match_out2877,
   input         match_out2878,
   input         match_out2879,
   input         match_out2880,
   input         match_out2881,
   input         match_out2882,
   input         match_out2883,
   input         match_out2884,
   input         match_out2885,
   input         match_out2886,
   input         match_out2887,
   input         match_out2888,
   input         match_out2889,
   input         match_out2890,
   input         match_out2891,
   input         match_out2892,
   input         match_out2893,
   input         match_out2894,
   input         match_out2895,
   input         match_out2896,
   input         match_out2897,
   input         match_out2898,
   input         match_out2899,
   input         match_out2900,
   input         match_out2901,
   input         match_out2902,
   input         match_out2903,
   input         match_out2904,
   input         match_out2905,
   input         match_out2906,
   input         match_out2907,
   input         match_out2908,
   input         match_out2909,
   input         match_out2910,
   input         match_out2911,
   input         match_out2912,
   input         match_out2913,
   input         match_out2914,
   input         match_out2915,
   input         match_out2916,
   input         match_out2917,
   input         match_out2918,
   input         match_out2919,
   input         match_out2920,
   input         match_out2921,
   input         match_out2922,
   input         match_out2923,
   input         match_out2924,
   input         match_out2925,
   input         match_out2926,
   input         match_out2927,
   input         match_out2928,
   input         match_out2929,
   input         match_out2930,
   input         match_out2931,
   input         match_out2932,
   input         match_out2933,
   input         match_out2934,
   input         match_out2935,
   input         match_out2936,
   input         match_out2937,
   input         match_out2938,
   input         match_out2939,
   input         match_out2940,
   input         match_out2941,
   input         match_out2942,
   input         match_out2943,
   input         match_out2944,
   input         match_out2945,
   input         match_out2946,
   input         match_out2947,
   input         match_out2948,
   input         match_out2949,
   input         match_out2950,
   input         match_out2951,
   input         match_out2952,
   input         match_out2953,
   input         match_out2954,
   input         match_out2955,
   input         match_out2956,
   input         match_out2957,
   input         match_out2958,
   input         match_out2959,
   input         match_out2960,
   input         match_out2961,
   input         match_out2962,
   input         match_out2963,
   input         match_out2964,
   input         match_out2965,
   input         match_out2966,
   input         match_out2967,
   input         match_out2968,
   input         match_out2969,
   input         match_out2970,
   input         match_out2971,
   input         match_out2972,
   input         match_out2973,
   input         match_out2974,
   input         match_out2975,
   input         match_out2976,
   input         match_out2977,
   input         match_out2978,
   input         match_out2979,
   input         match_out2980,
   input         match_out2981,
   input         match_out2982,
   input         match_out2983,
   input         match_out2984,
   input         match_out2985,
   input         match_out2986,
   input         match_out2987,
   input         match_out2988,
   input         match_out2989,
   input         match_out2990,
   input         match_out2991,
   input         match_out2992,
   input         match_out2993,
   input         match_out2994,
   input         match_out2995,
   input         match_out2996,
   input         match_out2997,
   input         match_out2998,
   input         match_out2999,
   input         match_out3000,
   input         match_out3001,
   input         match_out3002,
   input         match_out3003,
   input         match_out3004,
   input         match_out3005,
   input         match_out3006,
   input         match_out3007,
   input         match_out3008,
   input         match_out3009,
   input         match_out3010,
   input         match_out3011,
   input         match_out3012,
   input         match_out3013,
   input         match_out3014,
   input         match_out3015,
   input         match_out3016,
   input         match_out3017,
   input         match_out3018,
   input         match_out3019,
   input         match_out3020,
   input         match_out3021,
   input         match_out3022,
   input         match_out3023,
   input         match_out3024,
   input         match_out3025,
   input         match_out3026,
   input         match_out3027,
   input         match_out3028,
   input         match_out3029,
   input         match_out3030,
   input         match_out3031,
   input         match_out3032,
   input         match_out3033,
   input         match_out3034,
   input         match_out3035,
   input         match_out3036,
   input         match_out3037,
   input         match_out3038,
   input         match_out3039,
   input         match_out3040,
   input         match_out3041,
   input         match_out3042,
   input         match_out3043,
   input         match_out3044,
   input         match_out3045,
   input         match_out3046,
   input         match_out3047,
   input         match_out3048,
   input         match_out3049,
   input         match_out3050,
   input         match_out3051,
   input         match_out3052,
   input         match_out3053,
   input         match_out3054,
   input         match_out3055,
   input         match_out3056,
   input         match_out3057,
   input         match_out3058,
   input         match_out3059,
   input         match_out3060,
   input         match_out3061,
   input         match_out3062,
   input         match_out3063,
   input         match_out3064,
   input         match_out3065,
   input         match_out3066,
   input         match_out3067,
   input         match_out3068,
   input         match_out3069,
   input         match_out3070,
   input         match_out3071,
   input         match_out3072,
   input         match_out3073,
   input         match_out3074,
   input         match_out3075,
   input         match_out3076,
   input         match_out3077,
   input         match_out3078,
   input         match_out3079,
   input         match_out3080,
   input         match_out3081,
   input         match_out3082,
   input         match_out3083,
   input         match_out3084,
   input         match_out3085,
   input         match_out3086,
   input         match_out3087,
   input         match_out3088,
   input         match_out3089,
   input         match_out3090,
   input         match_out3091,
   input         match_out3092,
   input         match_out3093,
   input         match_out3094,
   input         match_out3095,
   input         match_out3096,
   input         match_out3097,
   input         match_out3098,
   input         match_out3099,
   input         match_out3100,
   input         match_out3101,
   input         match_out3102,
   input         match_out3103,
   input         match_out3104,
   input         match_out3105,
   input         match_out3106,
   input         match_out3107,
   input         match_out3108,
   input         match_out3109,
   input         match_out3110,
   input         match_out3111,
   input         match_out3112,
   input         match_out3113,
   input         match_out3114,
   input         match_out3115,
   input         match_out3116,
   input         match_out3117,
   input         match_out3118,
   input         match_out3119,
   input         match_out3120,
   input         match_out3121,
   input         match_out3122,
   input         match_out3123,
   input         match_out3124,
   input         match_out3125,
   input         match_out3126,
   input         match_out3127,
   input         match_out3128,
   input         match_out3129,
   input         match_out3130,
   input         match_out3131,
   input         match_out3132,
   input         match_out3133,
   input         match_out3134,
   input         match_out3135,
   input         match_out3136,
   input         match_out3137,
   input         match_out3138,
   input         match_out3139,
   input         match_out3140,
   input         match_out3141,
   input         match_out3142,
   input         match_out3143,
   input         match_out3144,
   input         match_out3145,
   input         match_out3146,
   input         match_out3147,
   input         match_out3148,
   input         match_out3149,
   input         match_out3150,
   input         match_out3151,
   input         match_out3152,
   input         match_out3153,
   input         match_out3154,
   input         match_out3155,
   input         match_out3156,
   input         match_out3157,
   input         match_out3158,
   input         match_out3159,
   input         match_out3160,
   input         match_out3161,
   input         match_out3162,
   input         match_out3163,
   input         match_out3164,
   input         match_out3165,
   input         match_out3166,
   input         match_out3167,
   input         match_out3168,
   input         match_out3169,
   input         match_out3170,
   input         match_out3171,
   input         match_out3172,
   input         match_out3173,
   input         match_out3174,
   input         match_out3175,
   input         match_out3176,
   input         match_out3177,
   input         match_out3178,
   input         match_out3179,
   input         match_out3180,
   input         match_out3181,
   input         match_out3182,
   input         match_out3183,
   input         match_out3184,
   input         match_out3185,
   input         match_out3186,
   input         match_out3187,
   input         match_out3188,
   input         match_out3189,
   input         match_out3190,
   input         match_out3191,
   input         match_out3192,
   input         match_out3193,
   input         match_out3194,
   input         match_out3195,
   input         match_out3196,
   input         match_out3197,
   input         match_out3198,
   input         match_out3199,
   input         match_out3200,
   input         match_out3201,
   input         match_out3202,
   input         match_out3203,
   input         match_out3204,
   input         match_out3205,
   input         match_out3206,
   input         match_out3207,
   input         match_out3208,
   input         match_out3209,
   input         match_out3210,
   input         match_out3211,
   input         match_out3212,
   input         match_out3213,
   input         match_out3214,
   input         match_out3215,
   input         match_out3216,
   input         match_out3217,
   input         match_out3218,
   input         match_out3219,
   input         match_out3220,
   input         match_out3221,
   input         match_out3222,
   input         match_out3223,
   input         match_out3224,
   input         match_out3225,
   input         match_out3226,
   input         match_out3227,
   input         match_out3228,
   input         match_out3229,
   input         match_out3230,
   input         match_out3231,
   input         match_out3232,
   input         match_out3233,
   input         match_out3234,
   input         match_out3235,
   input         match_out3236,
   input         match_out3237,
   input         match_out3238,
   input         match_out3239,
   input         match_out3240,
   input         match_out3241,
   input         match_out3242,
   input         match_out3243,
   input         match_out3244,
   input         match_out3245,
   input         match_out3246,
   input         match_out3247,
   input         match_out3248,
   input         match_out3249,
   input         match_out3250,
   input         match_out3251,
   input         match_out3252,
   input         match_out3253,
   input         match_out3254,
   input         match_out3255,
   input         match_out3256,
   input         match_out3257,
   input         match_out3258,
   input         match_out3259,
   input         match_out3260,
   input         match_out3261,
   input         match_out3262,
   input         match_out3263,
   input         match_out3264,
   input         match_out3265,
   input         match_out3266,
   input         match_out3267,
   input         match_out3268,
   input         match_out3269,
   input         match_out3270,
   input         match_out3271,
   input         match_out3272,
   input         match_out3273,
   input         match_out3274,
   input         match_out3275,
   input         match_out3276,
   input         match_out3277,
   input         match_out3278,
   input         match_out3279,
   input         match_out3280,
   input         match_out3281,
   input         match_out3282,
   input         match_out3283,
   input         match_out3284,
   input         match_out3285,
   input         match_out3286,
   input         match_out3287,
   input         match_out3288,
   input         match_out3289,
   input         match_out3290,
   input         match_out3291,
   input         match_out3292,
   input         match_out3293,
   input         match_out3294,
   input         match_out3295,
   input         match_out3296,
   input         match_out3297,
   input         match_out3298,
   input         match_out3299,
   input         match_out3300,
   input         match_out3301,
   input         match_out3302,
   input         match_out3303,
   input         match_out3304,
   input         match_out3305,
   input         match_out3306,
   input         match_out3307,
   input         match_out3308,
   input         match_out3309,
   input         match_out3310,
   input         match_out3311,
   input         match_out3312,
   input         match_out3313,
   input         match_out3314,
   input         match_out3315,
   input         match_out3316,
   input         match_out3317,
   input         match_out3318,
   input         match_out3319,
   input         match_out3320,
   input         match_out3321,
   input         match_out3322,
   input         match_out3323,
   input         match_out3324,
   input         match_out3325,
   input         match_out3326,
   input         match_out3327,
   input         match_out3328,
   input         match_out3329,
   input         match_out3330,
   input         match_out3331,
   input         match_out3332,
   input         match_out3333,
   input         match_out3334,
   input         match_out3335,
   input         match_out3336,
   input         match_out3337,
   input         match_out3338,
   input         match_out3339,
   input         match_out3340,
   input         match_out3341,
   input         match_out3342,
   input         match_out3343,
   input         match_out3344,
   input         match_out3345,
   input         match_out3346,
   input         match_out3347,
   input         match_out3348,
   input         match_out3349,
   input         match_out3350,
   input         match_out3351,
   input         match_out3352,
   input         match_out3353,
   input         match_out3354,
   input         match_out3355,
   input         match_out3356,
   input         match_out3357,
   input         match_out3358,
   input         match_out3359,
   input         match_out3360,
   input         match_out3361,
   input         match_out3362,
   input         match_out3363,
   input         match_out3364,
   input         match_out3365,
   input         match_out3366,
   input         match_out3367,
   input         match_out3368,
   input         match_out3369,
   input         match_out3370,
   input         match_out3371,
   input         match_out3372,
   input         match_out3373,
   input         match_out3374,
   input         match_out3375,
   input         match_out3376,
   input         match_out3377,
   input         match_out3378,
   input         match_out3379,
   input         match_out3380,
   input         match_out3381,
   input         match_out3382,
   input         match_out3383,
   input         match_out3384,
   input         match_out3385,
   input         match_out3386,
   input         match_out3387,
   input         match_out3388,
   input         match_out3389,
   input         match_out3390,
   input         match_out3391,
   input         match_out3392,
   input         match_out3393,
   input         match_out3394,
   input         match_out3395,
   input         match_out3396,
   input         match_out3397,
   input         match_out3398,
   input         match_out3399,
   input         match_out3400,
   input         match_out3401,
   input         match_out3402,
   input         match_out3403,
   input         match_out3404,
   input         match_out3405,
   input         match_out3406,
   input         match_out3407,
   input         match_out3408,
   input         match_out3409,
   input         match_out3410,
   input         match_out3411,
   input         match_out3412,
   input         match_out3413,
   input         match_out3414,
   input         match_out3415,
   input         match_out3416,
   input         match_out3417,
   input         match_out3418,
   input         match_out3419,
   input         match_out3420,
   input         match_out3421,
   input         match_out3422,
   input         match_out3423,
   input         match_out3424,
   input         match_out3425,
   input         match_out3426,
   input         match_out3427,
   input         match_out3428,
   input         match_out3429,
   input         match_out3430,
   input         match_out3431,
   input         match_out3432,
   input         match_out3433,
   input         match_out3434,
   input         match_out3435,
   input         match_out3436,
   input         match_out3437,
   input         match_out3438,
   input         match_out3439,
   input         match_out3440,
   input         match_out3441,
   input         match_out3442,
   input         match_out3443,
   input         match_out3444,
   input         match_out3445,
   input         match_out3446,
   input         match_out3447,
   input         match_out3448,
   input         match_out3449,
   input         match_out3450,
   input         match_out3451,
   input         match_out3452,
   input         match_out3453,
   input         match_out3454,
   input         match_out3455,
   input         match_out3456,
   input         match_out3457,
   input         match_out3458,
   input         match_out3459,
   input         match_out3460,
   input         match_out3461,
   input         match_out3462,
   input         match_out3463,
   input         match_out3464,
   input         match_out3465,
   input         match_out3466,
   input         match_out3467,
   input         match_out3468,
   input         match_out3469,
   input         match_out3470,
   input         match_out3471,
   input         match_out3472,
   input         match_out3473,
   input         match_out3474,
   input         match_out3475,
   input         match_out3476,
   input         match_out3477,
   input         match_out3478,
   input         match_out3479,
   input         match_out3480,
   input         match_out3481,
   input         match_out3482,
   input         match_out3483,
   input         match_out3484,
   input         match_out3485,
   input         match_out3486,
   input         match_out3487,
   input         match_out3488,
   input         match_out3489,
   input         match_out3490,
   input         match_out3491,
   input         match_out3492,
   input         match_out3493,
   input         match_out3494,
   input         match_out3495,
   input         match_out3496,
   input         match_out3497,
   input         match_out3498,
   input         match_out3499,
   input         match_out3500,
   input         match_out3501,
   input         match_out3502,
   input         match_out3503,
   input         match_out3504,
   input         match_out3505,
   input         match_out3506,
   input         match_out3507,
   input         match_out3508,
   input         match_out3509,
   input         match_out3510,
   input         match_out3511,
   input         match_out3512,
   input         match_out3513,
   input         match_out3514,
   input         match_out3515,
   input         match_out3516,
   input         match_out3517,
   input         match_out3518,
   input         match_out3519,
   input         match_out3520,
   input         match_out3521,
   input         match_out3522,
   input         match_out3523,
   input         match_out3524,
   input         match_out3525,
   input         match_out3526,
   input         match_out3527,
   input         match_out3528,
   input         match_out3529,
   input         match_out3530,
   input         match_out3531,
   input         match_out3532,
   input         match_out3533,
   input         match_out3534,
   input         match_out3535,
   input         match_out3536,
   input         match_out3537,
   input         match_out3538,
   input         match_out3539,
   input         match_out3540,
   input         match_out3541,
   input         match_out3542,
   input         match_out3543,
   input         match_out3544,
   input         match_out3545,
   input         match_out3546,
   input         match_out3547,
   input         match_out3548,
   input         match_out3549,
   input         match_out3550,
   input         match_out3551,
   input         match_out3552,
   input         match_out3553,
   input         match_out3554,
   input         match_out3555,
   input         match_out3556,
   input         match_out3557,
   input         match_out3558,
   input         match_out3559,
   input         match_out3560,
   input         match_out3561,
   input         match_out3562,
   input         match_out3563,
   input         match_out3564,
   input         match_out3565,
   input         match_out3566,
   input         match_out3567,
   input         match_out3568,
   input         match_out3569,
   input         match_out3570,
   input         match_out3571,
   input         match_out3572,
   input         match_out3573,
   input         match_out3574,
   input         match_out3575,
   input         match_out3576,
   input         match_out3577,
   input         match_out3578,
   input         match_out3579,
   input         match_out3580,
   input         match_out3581,
   input         match_out3582,
   input         match_out3583,
   input         match_out3584,
   input         match_out3585,
   input         match_out3586,
   input         match_out3587,
   input         match_out3588,
   input         match_out3589,
   input         match_out3590,
   input         match_out3591,
   input         match_out3592,
   input         match_out3593,
   input         match_out3594,
   input         match_out3595,
   input         match_out3596,
   input         match_out3597,
   input         match_out3598,
   input         match_out3599,
   input         match_out3600,
   input         match_out3601,
   input         match_out3602,
   input         match_out3603,
   input         match_out3604,
   input         match_out3605,
   input         match_out3606,
   input         match_out3607,
   input         match_out3608,
   input         match_out3609,
   input         match_out3610,
   input         match_out3611,
   input         match_out3612,
   input         match_out3613,
   input         match_out3614,
   input         match_out3615,
   input         match_out3616,
   input         match_out3617,
   input         match_out3618,
   input         match_out3619,
   input         match_out3620,
   input         match_out3621,
   input         match_out3622,
   input         match_out3623,
   input         match_out3624,
   input         match_out3625,
   input         match_out3626,
   input         match_out3627,
   input         match_out3628,
   input         match_out3629,
   input         match_out3630,
   input         match_out3631,
   input         match_out3632,
   input         match_out3633,
   input         match_out3634,
   input         match_out3635,
   input         match_out3636,
   input         match_out3637,
   input         match_out3638,
   input         match_out3639,
   input         match_out3640,
   input         match_out3641,
   input         match_out3642,
   input         match_out3643,
   input         match_out3644,
   input         match_out3645,
   input         match_out3646,
   input         match_out3647,
   input         match_out3648,
   input         match_out3649,
   input         match_out3650,
   input         match_out3651,
   input         match_out3652,
   input         match_out3653,
   input         match_out3654,
   input         match_out3655,
   input         match_out3656,
   input         match_out3657,
   input         match_out3658,
   input         match_out3659,
   input         match_out3660,
   input         match_out3661,
   input         match_out3662,
   input         match_out3663,
   input         match_out3664,
   input         match_out3665,
   input         match_out3666,
   input         match_out3667,
   input         match_out3668,
   input         match_out3669,
   input         match_out3670,
   input         match_out3671,
   input         match_out3672,
   input         match_out3673,
   input         match_out3674,
   input         match_out3675,
   input         match_out3676,
   input         match_out3677,
   input         match_out3678,
   input         match_out3679,
   input         match_out3680,
   input         match_out3681,
   input         match_out3682,
   input         match_out3683,
   input         match_out3684,
   input         match_out3685,
   input         match_out3686,
   input         match_out3687,
   input         match_out3688,
   input         match_out3689,
   input         match_out3690,
   input         match_out3691,
   input         match_out3692,
   input         match_out3693,
   input         match_out3694,
   input         match_out3695,
   input         match_out3696,
   input         match_out3697,
   input         match_out3698,
   input         match_out3699,
   input         match_out3700,
   input         match_out3701,
   input         match_out3702,
   input         match_out3703,
   input         match_out3704,
   input         match_out3705,
   input         match_out3706,
   input         match_out3707,
   input         match_out3708,
   input         match_out3709,
   input         match_out3710,
   input         match_out3711,
   input         match_out3712,
   input         match_out3713,
   input         match_out3714,
   input         match_out3715,
   input         match_out3716,
   input         match_out3717,
   input         match_out3718,
   input         match_out3719,
   input         match_out3720,
   input         match_out3721,
   input         match_out3722,
   input         match_out3723,
   input         match_out3724,
   input         match_out3725,
   input         match_out3726,
   input         match_out3727,
   input         match_out3728,
   input         match_out3729,
   input         match_out3730,
   input         match_out3731,
   input         match_out3732,
   input         match_out3733,
   input         match_out3734,
   input         match_out3735,
   input         match_out3736,
   input         match_out3737,
   input         match_out3738,
   input         match_out3739,
   input         match_out3740,
   input         match_out3741,
   input         match_out3742,
   input         match_out3743,
   input         match_out3744,
   input         match_out3745,
   input         match_out3746,
   input         match_out3747,
   input         match_out3748,
   input         match_out3749,
   input         match_out3750,
   input         match_out3751,
   input         match_out3752,
   input         match_out3753,
   input         match_out3754,
   input         match_out3755,
   input         match_out3756,
   input         match_out3757,
   input         match_out3758,
   input         match_out3759,
   input         match_out3760,
   input         match_out3761,
   input         match_out3762,
   input         match_out3763,
   input         match_out3764,
   input         match_out3765,
   input         match_out3766,
   input         match_out3767,
   input         match_out3768,
   input         match_out3769,
   input         match_out3770,
   input         match_out3771,
   input         match_out3772,
   input         match_out3773,
   input         match_out3774,
   input         match_out3775,
   input         match_out3776,
   input         match_out3777,
   input         match_out3778,
   input         match_out3779,
   input         match_out3780,
   input         match_out3781,
   input         match_out3782,
   input         match_out3783,
   input         match_out3784,
   input         match_out3785,
   input         match_out3786,
   input         match_out3787,
   input         match_out3788,
   input         match_out3789,
   input         match_out3790,
   input         match_out3791,
   input         match_out3792,
   input         match_out3793,
   input         match_out3794,
   input         match_out3795,
   input         match_out3796,
   input         match_out3797,
   input         match_out3798,
   input         match_out3799,
   input         match_out3800,
   input         match_out3801,
   input         match_out3802,
   input         match_out3803,
   input         match_out3804,
   input         match_out3805,
   input         match_out3806,
   input         match_out3807,
   input         match_out3808,
   input         match_out3809,
   input         match_out3810,
   input         match_out3811,
   input         match_out3812,
   input         match_out3813,
   input         match_out3814,
   input         match_out3815,
   input         match_out3816,
   input         match_out3817,
   input         match_out3818,
   input         match_out3819,
   input         match_out3820,
   input         match_out3821,
   input         match_out3822,
   input         match_out3823,
   input         match_out3824,
   input         match_out3825,
   input         match_out3826,
   input         match_out3827,
   input         match_out3828,
   input         match_out3829,
   input         match_out3830,
   input         match_out3831,
   input         match_out3832,
   input         match_out3833,
   input         match_out3834,
   input         match_out3835,
   input         match_out3836,
   input         match_out3837,
   input         match_out3838,
   input         match_out3839,
   input         match_out3840,
   input         match_out3841,
   input         match_out3842,
   input         match_out3843,
   input         match_out3844,
   input         match_out3845,
   input         match_out3846,
   input         match_out3847,
   input         match_out3848,
   input         match_out3849,
   input         match_out3850,
   input         match_out3851,
   input         match_out3852,
   input         match_out3853,
   input         match_out3854,
   input         match_out3855,
   input         match_out3856,
   input         match_out3857,
   input         match_out3858,
   input         match_out3859,
   input         match_out3860,
   input         match_out3861,
   input         match_out3862,
   input         match_out3863,
   input         match_out3864,
   input         match_out3865,
   input         match_out3866,
   input         match_out3867,
   input         match_out3868,
   input         match_out3869,
   input         match_out3870,
   input         match_out3871,
   input         match_out3872,
   input         match_out3873,
   input         match_out3874,
   input         match_out3875,
   input         match_out3876,
   input         match_out3877,
   input         match_out3878,
   input         match_out3879,
   input         match_out3880,
   input         match_out3881,
   input         match_out3882,
   input         match_out3883,
   input         match_out3884,
   input         match_out3885,
   input         match_out3886,
   input         match_out3887,
   input         match_out3888,
   input         match_out3889,
   input         match_out3890,
   input         match_out3891,
   input         match_out3892,
   input         match_out3893,
   input         match_out3894,
   input         match_out3895,
   input         match_out3896,
   input         match_out3897,
   input         match_out3898,
   input         match_out3899,
   input         match_out3900,
   input         match_out3901,
   input         match_out3902,
   input         match_out3903,
   input         match_out3904,
   input         match_out3905,
   input         match_out3906,
   input         match_out3907,
   input         match_out3908,
   input         match_out3909,
   input         match_out3910,
   input         match_out3911,
   input         match_out3912,
   input         match_out3913,
   input         match_out3914,
   input         match_out3915,
   input         match_out3916,
   input         match_out3917,
   input         match_out3918,
   input         match_out3919,
   input         match_out3920,
   input         match_out3921,
   input         match_out3922,
   input         match_out3923,
   input         match_out3924,
   input         match_out3925,
   input         match_out3926,
   input         match_out3927,
   input         match_out3928,
   input         match_out3929,
   input         match_out3930,
   input         match_out3931,
   input         match_out3932,
   input         match_out3933,
   input         match_out3934,
   input         match_out3935,
   input         match_out3936,
   input         match_out3937,
   input         match_out3938,
   input         match_out3939,
   input         match_out3940,
   input         match_out3941,
   input         match_out3942,
   input         match_out3943,
   input         match_out3944,
   input         match_out3945,
   input         match_out3946,
   input         match_out3947,
   input         match_out3948,
   input         match_out3949,
   input         match_out3950,
   input         match_out3951,
   input         match_out3952,
   input         match_out3953,
   input         match_out3954,
   input         match_out3955,
   input         match_out3956,
   input         match_out3957,
   input         match_out3958,
   input         match_out3959,
   input         match_out3960,
   input         match_out3961,
   input         match_out3962,
   input         match_out3963,
   input         match_out3964,
   input         match_out3965,
   input         match_out3966,
   input         match_out3967,
   input         match_out3968,
   input         match_out3969,
   input         match_out3970,
   input         match_out3971,
   input         match_out3972,
   input         match_out3973,
   input         match_out3974,
   input         match_out3975,
   input         match_out3976,
   input         match_out3977,
   input         match_out3978,
   input         match_out3979,
   input         match_out3980,
   input         match_out3981,
   input         match_out3982,
   input         match_out3983,
   input         match_out3984,
   input         match_out3985,
   input         match_out3986,
   input         match_out3987,
   input         match_out3988,
   input         match_out3989,
   input         match_out3990,
   input         match_out3991,
   input         match_out3992,
   input         match_out3993,
   input         match_out3994,
   input         match_out3995,
   input         match_out3996,
   input         match_out3997,
   input         match_out3998,
   input         match_out3999,
   input         match_out4000,
   input         match_out4001,
   input         match_out4002,
   input         match_out4003,
   input         match_out4004,
   input         match_out4005,
   input         match_out4006,
   input         match_out4007,
   input         match_out4008,
   input         match_out4009,
   input         match_out4010,
   input         match_out4011,
   input         match_out4012,
   input         match_out4013,
   input         match_out4014,
   input         match_out4015,
   input         match_out4016,
   input         match_out4017,
   input         match_out4018,
   input         match_out4019,
   input         match_out4020,
   input         match_out4021,
   input         match_out4022,
   input         match_out4023,
   input         match_out4024,
   input         match_out4025,
   input         match_out4026,
   input         match_out4027,
   input         match_out4028,
   input         match_out4029,
   input         match_out4030,
   input         match_out4031,
   input         match_out4032,
   input         match_out4033,
   input         match_out4034,
   input         match_out4035,
   input         match_out4036,
   input         match_out4037,
   input         match_out4038,
   input         match_out4039,
   input         match_out4040,
   input         match_out4041,
   input         match_out4042,
   input         match_out4043,
   input         match_out4044,
   input         match_out4045,
   input         match_out4046,
   input         match_out4047,
   input         match_out4048,
   input         match_out4049,
   input         match_out4050,
   input         match_out4051,
   input         match_out4052,
   input         match_out4053,
   input         match_out4054,
   input         match_out4055,
   input         match_out4056,
   input         match_out4057,
   input         match_out4058,
   input         match_out4059,
   input         match_out4060,
   input         match_out4061,
   input         match_out4062,
   input         match_out4063,
   input         match_out4064,
   input         match_out4065,
   input         match_out4066,
   input         match_out4067,
   input         match_out4068,
   input         match_out4069,
   input         match_out4070,
   input         match_out4071,
   input         match_out4072,
   input         match_out4073,
   input         match_out4074,
   input         match_out4075,
   input         match_out4076,
   input         match_out4077,
   input         match_out4078,
   input         match_out4079,
   input         match_out4080,
   input         match_out4081,
   input         match_out4082,
   input         match_out4083,
   input         match_out4084,
   input         match_out4085,
   input         match_out4086,
   input         match_out4087,
   input         match_out4088,
   input         match_out4089,
   input         match_out4090,
   input         match_out4091,
   input         match_out4092,
   input         match_out4093,
   input         match_out4094,
   input         match_out4095,
   output        cfg_en0,
   output        cfg_en1,
   output        cfg_en2,
   output        cfg_en3,
   output        cfg_en4,
   output        cfg_en5,
   output        cfg_en6,
   output        cfg_en7,
   output        cfg_en8,
   output        cfg_en9,
   output        cfg_en10,
   output        cfg_en11,
   output        cfg_en12,
   output        cfg_en13,
   output        cfg_en14,
   output        cfg_en15,
   output        cfg_en16,
   output        cfg_en17,
   output        cfg_en18,
   output        cfg_en19,
   output        cfg_en20,
   output        cfg_en21,
   output        cfg_en22,
   output        cfg_en23,
   output        cfg_en24,
   output        cfg_en25,
   output        cfg_en26,
   output        cfg_en27,
   output        cfg_en28,
   output        cfg_en29,
   output        cfg_en30,
   output        cfg_en31,
   output        cfg_en32,
   output        cfg_en33,
   output        cfg_en34,
   output        cfg_en35,
   output        cfg_en36,
   output        cfg_en37,
   output        cfg_en38,
   output        cfg_en39,
   output        cfg_en40,
   output        cfg_en41,
   output        cfg_en42,
   output        cfg_en43,
   output        cfg_en44,
   output        cfg_en45,
   output        cfg_en46,
   output        cfg_en47,
   output        cfg_en48,
   output        cfg_en49,
   output        cfg_en50,
   output        cfg_en51,
   output        cfg_en52,
   output        cfg_en53,
   output        cfg_en54,
   output        cfg_en55,
   output        cfg_en56,
   output        cfg_en57,
   output        cfg_en58,
   output        cfg_en59,
   output        cfg_en60,
   output        cfg_en61,
   output        cfg_en62,
   output        cfg_en63,
   output        cfg_en64,
   output        cfg_en65,
   output        cfg_en66,
   output        cfg_en67,
   output        cfg_en68,
   output        cfg_en69,
   output        cfg_en70,
   output        cfg_en71,
   output        cfg_en72,
   output        cfg_en73,
   output        cfg_en74,
   output        cfg_en75,
   output        cfg_en76,
   output        cfg_en77,
   output        cfg_en78,
   output        cfg_en79,
   output        cfg_en80,
   output        cfg_en81,
   output        cfg_en82,
   output        cfg_en83,
   output        cfg_en84,
   output        cfg_en85,
   output        cfg_en86,
   output        cfg_en87,
   output        cfg_en88,
   output        cfg_en89,
   output        cfg_en90,
   output        cfg_en91,
   output        cfg_en92,
   output        cfg_en93,
   output        cfg_en94,
   output        cfg_en95,
   output        cfg_en96,
   output        cfg_en97,
   output        cfg_en98,
   output        cfg_en99,
   output        cfg_en100,
   output        cfg_en101,
   output        cfg_en102,
   output        cfg_en103,
   output        cfg_en104,
   output        cfg_en105,
   output        cfg_en106,
   output        cfg_en107,
   output        cfg_en108,
   output        cfg_en109,
   output        cfg_en110,
   output        cfg_en111,
   output        cfg_en112,
   output        cfg_en113,
   output        cfg_en114,
   output        cfg_en115,
   output        cfg_en116,
   output        cfg_en117,
   output        cfg_en118,
   output        cfg_en119,
   output        cfg_en120,
   output        cfg_en121,
   output        cfg_en122,
   output        cfg_en123,
   output        cfg_en124,
   output        cfg_en125,
   output        cfg_en126,
   output        cfg_en127,
   output        cfg_en128,
   output        cfg_en129,
   output        cfg_en130,
   output        cfg_en131,
   output        cfg_en132,
   output        cfg_en133,
   output        cfg_en134,
   output        cfg_en135,
   output        cfg_en136,
   output        cfg_en137,
   output        cfg_en138,
   output        cfg_en139,
   output        cfg_en140,
   output        cfg_en141,
   output        cfg_en142,
   output        cfg_en143,
   output        cfg_en144,
   output        cfg_en145,
   output        cfg_en146,
   output        cfg_en147,
   output        cfg_en148,
   output        cfg_en149,
   output        cfg_en150,
   output        cfg_en151,
   output        cfg_en152,
   output        cfg_en153,
   output        cfg_en154,
   output        cfg_en155,
   output        cfg_en156,
   output        cfg_en157,
   output        cfg_en158,
   output        cfg_en159,
   output        cfg_en160,
   output        cfg_en161,
   output        cfg_en162,
   output        cfg_en163,
   output        cfg_en164,
   output        cfg_en165,
   output        cfg_en166,
   output        cfg_en167,
   output        cfg_en168,
   output        cfg_en169,
   output        cfg_en170,
   output        cfg_en171,
   output        cfg_en172,
   output        cfg_en173,
   output        cfg_en174,
   output        cfg_en175,
   output        cfg_en176,
   output        cfg_en177,
   output        cfg_en178,
   output        cfg_en179,
   output        cfg_en180,
   output        cfg_en181,
   output        cfg_en182,
   output        cfg_en183,
   output        cfg_en184,
   output        cfg_en185,
   output        cfg_en186,
   output        cfg_en187,
   output        cfg_en188,
   output        cfg_en189,
   output        cfg_en190,
   output        cfg_en191,
   output        cfg_en192,
   output        cfg_en193,
   output        cfg_en194,
   output        cfg_en195,
   output        cfg_en196,
   output        cfg_en197,
   output        cfg_en198,
   output        cfg_en199,
   output        cfg_en200,
   output        cfg_en201,
   output        cfg_en202,
   output        cfg_en203,
   output        cfg_en204,
   output        cfg_en205,
   output        cfg_en206,
   output        cfg_en207,
   output        cfg_en208,
   output        cfg_en209,
   output        cfg_en210,
   output        cfg_en211,
   output        cfg_en212,
   output        cfg_en213,
   output        cfg_en214,
   output        cfg_en215,
   output        cfg_en216,
   output        cfg_en217,
   output        cfg_en218,
   output        cfg_en219,
   output        cfg_en220,
   output        cfg_en221,
   output        cfg_en222,
   output        cfg_en223,
   output        cfg_en224,
   output        cfg_en225,
   output        cfg_en226,
   output        cfg_en227,
   output        cfg_en228,
   output        cfg_en229,
   output        cfg_en230,
   output        cfg_en231,
   output        cfg_en232,
   output        cfg_en233,
   output        cfg_en234,
   output        cfg_en235,
   output        cfg_en236,
   output        cfg_en237,
   output        cfg_en238,
   output        cfg_en239,
   output        cfg_en240,
   output        cfg_en241,
   output        cfg_en242,
   output        cfg_en243,
   output        cfg_en244,
   output        cfg_en245,
   output        cfg_en246,
   output        cfg_en247,
   output        cfg_en248,
   output        cfg_en249,
   output        cfg_en250,
   output        cfg_en251,
   output        cfg_en252,
   output        cfg_en253,
   output        cfg_en254,
   output        cfg_en255,
   output        cfg_en256,
   output        cfg_en257,
   output        cfg_en258,
   output        cfg_en259,
   output        cfg_en260,
   output        cfg_en261,
   output        cfg_en262,
   output        cfg_en263,
   output        cfg_en264,
   output        cfg_en265,
   output        cfg_en266,
   output        cfg_en267,
   output        cfg_en268,
   output        cfg_en269,
   output        cfg_en270,
   output        cfg_en271,
   output        cfg_en272,
   output        cfg_en273,
   output        cfg_en274,
   output        cfg_en275,
   output        cfg_en276,
   output        cfg_en277,
   output        cfg_en278,
   output        cfg_en279,
   output        cfg_en280,
   output        cfg_en281,
   output        cfg_en282,
   output        cfg_en283,
   output        cfg_en284,
   output        cfg_en285,
   output        cfg_en286,
   output        cfg_en287,
   output        cfg_en288,
   output        cfg_en289,
   output        cfg_en290,
   output        cfg_en291,
   output        cfg_en292,
   output        cfg_en293,
   output        cfg_en294,
   output        cfg_en295,
   output        cfg_en296,
   output        cfg_en297,
   output        cfg_en298,
   output        cfg_en299,
   output        cfg_en300,
   output        cfg_en301,
   output        cfg_en302,
   output        cfg_en303,
   output        cfg_en304,
   output        cfg_en305,
   output        cfg_en306,
   output        cfg_en307,
   output        cfg_en308,
   output        cfg_en309,
   output        cfg_en310,
   output        cfg_en311,
   output        cfg_en312,
   output        cfg_en313,
   output        cfg_en314,
   output        cfg_en315,
   output        cfg_en316,
   output        cfg_en317,
   output        cfg_en318,
   output        cfg_en319,
   output        cfg_en320,
   output        cfg_en321,
   output        cfg_en322,
   output        cfg_en323,
   output        cfg_en324,
   output        cfg_en325,
   output        cfg_en326,
   output        cfg_en327,
   output        cfg_en328,
   output        cfg_en329,
   output        cfg_en330,
   output        cfg_en331,
   output        cfg_en332,
   output        cfg_en333,
   output        cfg_en334,
   output        cfg_en335,
   output        cfg_en336,
   output        cfg_en337,
   output        cfg_en338,
   output        cfg_en339,
   output        cfg_en340,
   output        cfg_en341,
   output        cfg_en342,
   output        cfg_en343,
   output        cfg_en344,
   output        cfg_en345,
   output        cfg_en346,
   output        cfg_en347,
   output        cfg_en348,
   output        cfg_en349,
   output        cfg_en350,
   output        cfg_en351,
   output        cfg_en352,
   output        cfg_en353,
   output        cfg_en354,
   output        cfg_en355,
   output        cfg_en356,
   output        cfg_en357,
   output        cfg_en358,
   output        cfg_en359,
   output        cfg_en360,
   output        cfg_en361,
   output        cfg_en362,
   output        cfg_en363,
   output        cfg_en364,
   output        cfg_en365,
   output        cfg_en366,
   output        cfg_en367,
   output        cfg_en368,
   output        cfg_en369,
   output        cfg_en370,
   output        cfg_en371,
   output        cfg_en372,
   output        cfg_en373,
   output        cfg_en374,
   output        cfg_en375,
   output        cfg_en376,
   output        cfg_en377,
   output        cfg_en378,
   output        cfg_en379,
   output        cfg_en380,
   output        cfg_en381,
   output        cfg_en382,
   output        cfg_en383,
   output        cfg_en384,
   output        cfg_en385,
   output        cfg_en386,
   output        cfg_en387,
   output        cfg_en388,
   output        cfg_en389,
   output        cfg_en390,
   output        cfg_en391,
   output        cfg_en392,
   output        cfg_en393,
   output        cfg_en394,
   output        cfg_en395,
   output        cfg_en396,
   output        cfg_en397,
   output        cfg_en398,
   output        cfg_en399,
   output        cfg_en400,
   output        cfg_en401,
   output        cfg_en402,
   output        cfg_en403,
   output        cfg_en404,
   output        cfg_en405,
   output        cfg_en406,
   output        cfg_en407,
   output        cfg_en408,
   output        cfg_en409,
   output        cfg_en410,
   output        cfg_en411,
   output        cfg_en412,
   output        cfg_en413,
   output        cfg_en414,
   output        cfg_en415,
   output        cfg_en416,
   output        cfg_en417,
   output        cfg_en418,
   output        cfg_en419,
   output        cfg_en420,
   output        cfg_en421,
   output        cfg_en422,
   output        cfg_en423,
   output        cfg_en424,
   output        cfg_en425,
   output        cfg_en426,
   output        cfg_en427,
   output        cfg_en428,
   output        cfg_en429,
   output        cfg_en430,
   output        cfg_en431,
   output        cfg_en432,
   output        cfg_en433,
   output        cfg_en434,
   output        cfg_en435,
   output        cfg_en436,
   output        cfg_en437,
   output        cfg_en438,
   output        cfg_en439,
   output        cfg_en440,
   output        cfg_en441,
   output        cfg_en442,
   output        cfg_en443,
   output        cfg_en444,
   output        cfg_en445,
   output        cfg_en446,
   output        cfg_en447,
   output        cfg_en448,
   output        cfg_en449,
   output        cfg_en450,
   output        cfg_en451,
   output        cfg_en452,
   output        cfg_en453,
   output        cfg_en454,
   output        cfg_en455,
   output        cfg_en456,
   output        cfg_en457,
   output        cfg_en458,
   output        cfg_en459,
   output        cfg_en460,
   output        cfg_en461,
   output        cfg_en462,
   output        cfg_en463,
   output        cfg_en464,
   output        cfg_en465,
   output        cfg_en466,
   output        cfg_en467,
   output        cfg_en468,
   output        cfg_en469,
   output        cfg_en470,
   output        cfg_en471,
   output        cfg_en472,
   output        cfg_en473,
   output        cfg_en474,
   output        cfg_en475,
   output        cfg_en476,
   output        cfg_en477,
   output        cfg_en478,
   output        cfg_en479,
   output        cfg_en480,
   output        cfg_en481,
   output        cfg_en482,
   output        cfg_en483,
   output        cfg_en484,
   output        cfg_en485,
   output        cfg_en486,
   output        cfg_en487,
   output        cfg_en488,
   output        cfg_en489,
   output        cfg_en490,
   output        cfg_en491,
   output        cfg_en492,
   output        cfg_en493,
   output        cfg_en494,
   output        cfg_en495,
   output        cfg_en496,
   output        cfg_en497,
   output        cfg_en498,
   output        cfg_en499,
   output        cfg_en500,
   output        cfg_en501,
   output        cfg_en502,
   output        cfg_en503,
   output        cfg_en504,
   output        cfg_en505,
   output        cfg_en506,
   output        cfg_en507,
   output        cfg_en508,
   output        cfg_en509,
   output        cfg_en510,
   output        cfg_en511,
   output        cfg_en512,
   output        cfg_en513,
   output        cfg_en514,
   output        cfg_en515,
   output        cfg_en516,
   output        cfg_en517,
   output        cfg_en518,
   output        cfg_en519,
   output        cfg_en520,
   output        cfg_en521,
   output        cfg_en522,
   output        cfg_en523,
   output        cfg_en524,
   output        cfg_en525,
   output        cfg_en526,
   output        cfg_en527,
   output        cfg_en528,
   output        cfg_en529,
   output        cfg_en530,
   output        cfg_en531,
   output        cfg_en532,
   output        cfg_en533,
   output        cfg_en534,
   output        cfg_en535,
   output        cfg_en536,
   output        cfg_en537,
   output        cfg_en538,
   output        cfg_en539,
   output        cfg_en540,
   output        cfg_en541,
   output        cfg_en542,
   output        cfg_en543,
   output        cfg_en544,
   output        cfg_en545,
   output        cfg_en546,
   output        cfg_en547,
   output        cfg_en548,
   output        cfg_en549,
   output        cfg_en550,
   output        cfg_en551,
   output        cfg_en552,
   output        cfg_en553,
   output        cfg_en554,
   output        cfg_en555,
   output        cfg_en556,
   output        cfg_en557,
   output        cfg_en558,
   output        cfg_en559,
   output        cfg_en560,
   output        cfg_en561,
   output        cfg_en562,
   output        cfg_en563,
   output        cfg_en564,
   output        cfg_en565,
   output        cfg_en566,
   output        cfg_en567,
   output        cfg_en568,
   output        cfg_en569,
   output        cfg_en570,
   output        cfg_en571,
   output        cfg_en572,
   output        cfg_en573,
   output        cfg_en574,
   output        cfg_en575,
   output        cfg_en576,
   output        cfg_en577,
   output        cfg_en578,
   output        cfg_en579,
   output        cfg_en580,
   output        cfg_en581,
   output        cfg_en582,
   output        cfg_en583,
   output        cfg_en584,
   output        cfg_en585,
   output        cfg_en586,
   output        cfg_en587,
   output        cfg_en588,
   output        cfg_en589,
   output        cfg_en590,
   output        cfg_en591,
   output        cfg_en592,
   output        cfg_en593,
   output        cfg_en594,
   output        cfg_en595,
   output        cfg_en596,
   output        cfg_en597,
   output        cfg_en598,
   output        cfg_en599,
   output        cfg_en600,
   output        cfg_en601,
   output        cfg_en602,
   output        cfg_en603,
   output        cfg_en604,
   output        cfg_en605,
   output        cfg_en606,
   output        cfg_en607,
   output        cfg_en608,
   output        cfg_en609,
   output        cfg_en610,
   output        cfg_en611,
   output        cfg_en612,
   output        cfg_en613,
   output        cfg_en614,
   output        cfg_en615,
   output        cfg_en616,
   output        cfg_en617,
   output        cfg_en618,
   output        cfg_en619,
   output        cfg_en620,
   output        cfg_en621,
   output        cfg_en622,
   output        cfg_en623,
   output        cfg_en624,
   output        cfg_en625,
   output        cfg_en626,
   output        cfg_en627,
   output        cfg_en628,
   output        cfg_en629,
   output        cfg_en630,
   output        cfg_en631,
   output        cfg_en632,
   output        cfg_en633,
   output        cfg_en634,
   output        cfg_en635,
   output        cfg_en636,
   output        cfg_en637,
   output        cfg_en638,
   output        cfg_en639,
   output        cfg_en640,
   output        cfg_en641,
   output        cfg_en642,
   output        cfg_en643,
   output        cfg_en644,
   output        cfg_en645,
   output        cfg_en646,
   output        cfg_en647,
   output        cfg_en648,
   output        cfg_en649,
   output        cfg_en650,
   output        cfg_en651,
   output        cfg_en652,
   output        cfg_en653,
   output        cfg_en654,
   output        cfg_en655,
   output        cfg_en656,
   output        cfg_en657,
   output        cfg_en658,
   output        cfg_en659,
   output        cfg_en660,
   output        cfg_en661,
   output        cfg_en662,
   output        cfg_en663,
   output        cfg_en664,
   output        cfg_en665,
   output        cfg_en666,
   output        cfg_en667,
   output        cfg_en668,
   output        cfg_en669,
   output        cfg_en670,
   output        cfg_en671,
   output        cfg_en672,
   output        cfg_en673,
   output        cfg_en674,
   output        cfg_en675,
   output        cfg_en676,
   output        cfg_en677,
   output        cfg_en678,
   output        cfg_en679,
   output        cfg_en680,
   output        cfg_en681,
   output        cfg_en682,
   output        cfg_en683,
   output        cfg_en684,
   output        cfg_en685,
   output        cfg_en686,
   output        cfg_en687,
   output        cfg_en688,
   output        cfg_en689,
   output        cfg_en690,
   output        cfg_en691,
   output        cfg_en692,
   output        cfg_en693,
   output        cfg_en694,
   output        cfg_en695,
   output        cfg_en696,
   output        cfg_en697,
   output        cfg_en698,
   output        cfg_en699,
   output        cfg_en700,
   output        cfg_en701,
   output        cfg_en702,
   output        cfg_en703,
   output        cfg_en704,
   output        cfg_en705,
   output        cfg_en706,
   output        cfg_en707,
   output        cfg_en708,
   output        cfg_en709,
   output        cfg_en710,
   output        cfg_en711,
   output        cfg_en712,
   output        cfg_en713,
   output        cfg_en714,
   output        cfg_en715,
   output        cfg_en716,
   output        cfg_en717,
   output        cfg_en718,
   output        cfg_en719,
   output        cfg_en720,
   output        cfg_en721,
   output        cfg_en722,
   output        cfg_en723,
   output        cfg_en724,
   output        cfg_en725,
   output        cfg_en726,
   output        cfg_en727,
   output        cfg_en728,
   output        cfg_en729,
   output        cfg_en730,
   output        cfg_en731,
   output        cfg_en732,
   output        cfg_en733,
   output        cfg_en734,
   output        cfg_en735,
   output        cfg_en736,
   output        cfg_en737,
   output        cfg_en738,
   output        cfg_en739,
   output        cfg_en740,
   output        cfg_en741,
   output        cfg_en742,
   output        cfg_en743,
   output        cfg_en744,
   output        cfg_en745,
   output        cfg_en746,
   output        cfg_en747,
   output        cfg_en748,
   output        cfg_en749,
   output        cfg_en750,
   output        cfg_en751,
   output        cfg_en752,
   output        cfg_en753,
   output        cfg_en754,
   output        cfg_en755,
   output        cfg_en756,
   output        cfg_en757,
   output        cfg_en758,
   output        cfg_en759,
   output        cfg_en760,
   output        cfg_en761,
   output        cfg_en762,
   output        cfg_en763,
   output        cfg_en764,
   output        cfg_en765,
   output        cfg_en766,
   output        cfg_en767,
   output        cfg_en768,
   output        cfg_en769,
   output        cfg_en770,
   output        cfg_en771,
   output        cfg_en772,
   output        cfg_en773,
   output        cfg_en774,
   output        cfg_en775,
   output        cfg_en776,
   output        cfg_en777,
   output        cfg_en778,
   output        cfg_en779,
   output        cfg_en780,
   output        cfg_en781,
   output        cfg_en782,
   output        cfg_en783,
   output        cfg_en784,
   output        cfg_en785,
   output        cfg_en786,
   output        cfg_en787,
   output        cfg_en788,
   output        cfg_en789,
   output        cfg_en790,
   output        cfg_en791,
   output        cfg_en792,
   output        cfg_en793,
   output        cfg_en794,
   output        cfg_en795,
   output        cfg_en796,
   output        cfg_en797,
   output        cfg_en798,
   output        cfg_en799,
   output        cfg_en800,
   output        cfg_en801,
   output        cfg_en802,
   output        cfg_en803,
   output        cfg_en804,
   output        cfg_en805,
   output        cfg_en806,
   output        cfg_en807,
   output        cfg_en808,
   output        cfg_en809,
   output        cfg_en810,
   output        cfg_en811,
   output        cfg_en812,
   output        cfg_en813,
   output        cfg_en814,
   output        cfg_en815,
   output        cfg_en816,
   output        cfg_en817,
   output        cfg_en818,
   output        cfg_en819,
   output        cfg_en820,
   output        cfg_en821,
   output        cfg_en822,
   output        cfg_en823,
   output        cfg_en824,
   output        cfg_en825,
   output        cfg_en826,
   output        cfg_en827,
   output        cfg_en828,
   output        cfg_en829,
   output        cfg_en830,
   output        cfg_en831,
   output        cfg_en832,
   output        cfg_en833,
   output        cfg_en834,
   output        cfg_en835,
   output        cfg_en836,
   output        cfg_en837,
   output        cfg_en838,
   output        cfg_en839,
   output        cfg_en840,
   output        cfg_en841,
   output        cfg_en842,
   output        cfg_en843,
   output        cfg_en844,
   output        cfg_en845,
   output        cfg_en846,
   output        cfg_en847,
   output        cfg_en848,
   output        cfg_en849,
   output        cfg_en850,
   output        cfg_en851,
   output        cfg_en852,
   output        cfg_en853,
   output        cfg_en854,
   output        cfg_en855,
   output        cfg_en856,
   output        cfg_en857,
   output        cfg_en858,
   output        cfg_en859,
   output        cfg_en860,
   output        cfg_en861,
   output        cfg_en862,
   output        cfg_en863,
   output        cfg_en864,
   output        cfg_en865,
   output        cfg_en866,
   output        cfg_en867,
   output        cfg_en868,
   output        cfg_en869,
   output        cfg_en870,
   output        cfg_en871,
   output        cfg_en872,
   output        cfg_en873,
   output        cfg_en874,
   output        cfg_en875,
   output        cfg_en876,
   output        cfg_en877,
   output        cfg_en878,
   output        cfg_en879,
   output        cfg_en880,
   output        cfg_en881,
   output        cfg_en882,
   output        cfg_en883,
   output        cfg_en884,
   output        cfg_en885,
   output        cfg_en886,
   output        cfg_en887,
   output        cfg_en888,
   output        cfg_en889,
   output        cfg_en890,
   output        cfg_en891,
   output        cfg_en892,
   output        cfg_en893,
   output        cfg_en894,
   output        cfg_en895,
   output        cfg_en896,
   output        cfg_en897,
   output        cfg_en898,
   output        cfg_en899,
   output        cfg_en900,
   output        cfg_en901,
   output        cfg_en902,
   output        cfg_en903,
   output        cfg_en904,
   output        cfg_en905,
   output        cfg_en906,
   output        cfg_en907,
   output        cfg_en908,
   output        cfg_en909,
   output        cfg_en910,
   output        cfg_en911,
   output        cfg_en912,
   output        cfg_en913,
   output        cfg_en914,
   output        cfg_en915,
   output        cfg_en916,
   output        cfg_en917,
   output        cfg_en918,
   output        cfg_en919,
   output        cfg_en920,
   output        cfg_en921,
   output        cfg_en922,
   output        cfg_en923,
   output        cfg_en924,
   output        cfg_en925,
   output        cfg_en926,
   output        cfg_en927,
   output        cfg_en928,
   output        cfg_en929,
   output        cfg_en930,
   output        cfg_en931,
   output        cfg_en932,
   output        cfg_en933,
   output        cfg_en934,
   output        cfg_en935,
   output        cfg_en936,
   output        cfg_en937,
   output        cfg_en938,
   output        cfg_en939,
   output        cfg_en940,
   output        cfg_en941,
   output        cfg_en942,
   output        cfg_en943,
   output        cfg_en944,
   output        cfg_en945,
   output        cfg_en946,
   output        cfg_en947,
   output        cfg_en948,
   output        cfg_en949,
   output        cfg_en950,
   output        cfg_en951,
   output        cfg_en952,
   output        cfg_en953,
   output        cfg_en954,
   output        cfg_en955,
   output        cfg_en956,
   output        cfg_en957,
   output        cfg_en958,
   output        cfg_en959,
   output        cfg_en960,
   output        cfg_en961,
   output        cfg_en962,
   output        cfg_en963,
   output        cfg_en964,
   output        cfg_en965,
   output        cfg_en966,
   output        cfg_en967,
   output        cfg_en968,
   output        cfg_en969,
   output        cfg_en970,
   output        cfg_en971,
   output        cfg_en972,
   output        cfg_en973,
   output        cfg_en974,
   output        cfg_en975,
   output        cfg_en976,
   output        cfg_en977,
   output        cfg_en978,
   output        cfg_en979,
   output        cfg_en980,
   output        cfg_en981,
   output        cfg_en982,
   output        cfg_en983,
   output        cfg_en984,
   output        cfg_en985,
   output        cfg_en986,
   output        cfg_en987,
   output        cfg_en988,
   output        cfg_en989,
   output        cfg_en990,
   output        cfg_en991,
   output        cfg_en992,
   output        cfg_en993,
   output        cfg_en994,
   output        cfg_en995,
   output        cfg_en996,
   output        cfg_en997,
   output        cfg_en998,
   output        cfg_en999,
   output        cfg_en1000,
   output        cfg_en1001,
   output        cfg_en1002,
   output        cfg_en1003,
   output        cfg_en1004,
   output        cfg_en1005,
   output        cfg_en1006,
   output        cfg_en1007,
   output        cfg_en1008,
   output        cfg_en1009,
   output        cfg_en1010,
   output        cfg_en1011,
   output        cfg_en1012,
   output        cfg_en1013,
   output        cfg_en1014,
   output        cfg_en1015,
   output        cfg_en1016,
   output        cfg_en1017,
   output        cfg_en1018,
   output        cfg_en1019,
   output        cfg_en1020,
   output        cfg_en1021,
   output        cfg_en1022,
   output        cfg_en1023,
   output        cfg_en1024,
   output        cfg_en1025,
   output        cfg_en1026,
   output        cfg_en1027,
   output        cfg_en1028,
   output        cfg_en1029,
   output        cfg_en1030,
   output        cfg_en1031,
   output        cfg_en1032,
   output        cfg_en1033,
   output        cfg_en1034,
   output        cfg_en1035,
   output        cfg_en1036,
   output        cfg_en1037,
   output        cfg_en1038,
   output        cfg_en1039,
   output        cfg_en1040,
   output        cfg_en1041,
   output        cfg_en1042,
   output        cfg_en1043,
   output        cfg_en1044,
   output        cfg_en1045,
   output        cfg_en1046,
   output        cfg_en1047,
   output        cfg_en1048,
   output        cfg_en1049,
   output        cfg_en1050,
   output        cfg_en1051,
   output        cfg_en1052,
   output        cfg_en1053,
   output        cfg_en1054,
   output        cfg_en1055,
   output        cfg_en1056,
   output        cfg_en1057,
   output        cfg_en1058,
   output        cfg_en1059,
   output        cfg_en1060,
   output        cfg_en1061,
   output        cfg_en1062,
   output        cfg_en1063,
   output        cfg_en1064,
   output        cfg_en1065,
   output        cfg_en1066,
   output        cfg_en1067,
   output        cfg_en1068,
   output        cfg_en1069,
   output        cfg_en1070,
   output        cfg_en1071,
   output        cfg_en1072,
   output        cfg_en1073,
   output        cfg_en1074,
   output        cfg_en1075,
   output        cfg_en1076,
   output        cfg_en1077,
   output        cfg_en1078,
   output        cfg_en1079,
   output        cfg_en1080,
   output        cfg_en1081,
   output        cfg_en1082,
   output        cfg_en1083,
   output        cfg_en1084,
   output        cfg_en1085,
   output        cfg_en1086,
   output        cfg_en1087,
   output        cfg_en1088,
   output        cfg_en1089,
   output        cfg_en1090,
   output        cfg_en1091,
   output        cfg_en1092,
   output        cfg_en1093,
   output        cfg_en1094,
   output        cfg_en1095,
   output        cfg_en1096,
   output        cfg_en1097,
   output        cfg_en1098,
   output        cfg_en1099,
   output        cfg_en1100,
   output        cfg_en1101,
   output        cfg_en1102,
   output        cfg_en1103,
   output        cfg_en1104,
   output        cfg_en1105,
   output        cfg_en1106,
   output        cfg_en1107,
   output        cfg_en1108,
   output        cfg_en1109,
   output        cfg_en1110,
   output        cfg_en1111,
   output        cfg_en1112,
   output        cfg_en1113,
   output        cfg_en1114,
   output        cfg_en1115,
   output        cfg_en1116,
   output        cfg_en1117,
   output        cfg_en1118,
   output        cfg_en1119,
   output        cfg_en1120,
   output        cfg_en1121,
   output        cfg_en1122,
   output        cfg_en1123,
   output        cfg_en1124,
   output        cfg_en1125,
   output        cfg_en1126,
   output        cfg_en1127,
   output        cfg_en1128,
   output        cfg_en1129,
   output        cfg_en1130,
   output        cfg_en1131,
   output        cfg_en1132,
   output        cfg_en1133,
   output        cfg_en1134,
   output        cfg_en1135,
   output        cfg_en1136,
   output        cfg_en1137,
   output        cfg_en1138,
   output        cfg_en1139,
   output        cfg_en1140,
   output        cfg_en1141,
   output        cfg_en1142,
   output        cfg_en1143,
   output        cfg_en1144,
   output        cfg_en1145,
   output        cfg_en1146,
   output        cfg_en1147,
   output        cfg_en1148,
   output        cfg_en1149,
   output        cfg_en1150,
   output        cfg_en1151,
   output        cfg_en1152,
   output        cfg_en1153,
   output        cfg_en1154,
   output        cfg_en1155,
   output        cfg_en1156,
   output        cfg_en1157,
   output        cfg_en1158,
   output        cfg_en1159,
   output        cfg_en1160,
   output        cfg_en1161,
   output        cfg_en1162,
   output        cfg_en1163,
   output        cfg_en1164,
   output        cfg_en1165,
   output        cfg_en1166,
   output        cfg_en1167,
   output        cfg_en1168,
   output        cfg_en1169,
   output        cfg_en1170,
   output        cfg_en1171,
   output        cfg_en1172,
   output        cfg_en1173,
   output        cfg_en1174,
   output        cfg_en1175,
   output        cfg_en1176,
   output        cfg_en1177,
   output        cfg_en1178,
   output        cfg_en1179,
   output        cfg_en1180,
   output        cfg_en1181,
   output        cfg_en1182,
   output        cfg_en1183,
   output        cfg_en1184,
   output        cfg_en1185,
   output        cfg_en1186,
   output        cfg_en1187,
   output        cfg_en1188,
   output        cfg_en1189,
   output        cfg_en1190,
   output        cfg_en1191,
   output        cfg_en1192,
   output        cfg_en1193,
   output        cfg_en1194,
   output        cfg_en1195,
   output        cfg_en1196,
   output        cfg_en1197,
   output        cfg_en1198,
   output        cfg_en1199,
   output        cfg_en1200,
   output        cfg_en1201,
   output        cfg_en1202,
   output        cfg_en1203,
   output        cfg_en1204,
   output        cfg_en1205,
   output        cfg_en1206,
   output        cfg_en1207,
   output        cfg_en1208,
   output        cfg_en1209,
   output        cfg_en1210,
   output        cfg_en1211,
   output        cfg_en1212,
   output        cfg_en1213,
   output        cfg_en1214,
   output        cfg_en1215,
   output        cfg_en1216,
   output        cfg_en1217,
   output        cfg_en1218,
   output        cfg_en1219,
   output        cfg_en1220,
   output        cfg_en1221,
   output        cfg_en1222,
   output        cfg_en1223,
   output        cfg_en1224,
   output        cfg_en1225,
   output        cfg_en1226,
   output        cfg_en1227,
   output        cfg_en1228,
   output        cfg_en1229,
   output        cfg_en1230,
   output        cfg_en1231,
   output        cfg_en1232,
   output        cfg_en1233,
   output        cfg_en1234,
   output        cfg_en1235,
   output        cfg_en1236,
   output        cfg_en1237,
   output        cfg_en1238,
   output        cfg_en1239,
   output        cfg_en1240,
   output        cfg_en1241,
   output        cfg_en1242,
   output        cfg_en1243,
   output        cfg_en1244,
   output        cfg_en1245,
   output        cfg_en1246,
   output        cfg_en1247,
   output        cfg_en1248,
   output        cfg_en1249,
   output        cfg_en1250,
   output        cfg_en1251,
   output        cfg_en1252,
   output        cfg_en1253,
   output        cfg_en1254,
   output        cfg_en1255,
   output        cfg_en1256,
   output        cfg_en1257,
   output        cfg_en1258,
   output        cfg_en1259,
   output        cfg_en1260,
   output        cfg_en1261,
   output        cfg_en1262,
   output        cfg_en1263,
   output        cfg_en1264,
   output        cfg_en1265,
   output        cfg_en1266,
   output        cfg_en1267,
   output        cfg_en1268,
   output        cfg_en1269,
   output        cfg_en1270,
   output        cfg_en1271,
   output        cfg_en1272,
   output        cfg_en1273,
   output        cfg_en1274,
   output        cfg_en1275,
   output        cfg_en1276,
   output        cfg_en1277,
   output        cfg_en1278,
   output        cfg_en1279,
   output        cfg_en1280,
   output        cfg_en1281,
   output        cfg_en1282,
   output        cfg_en1283,
   output        cfg_en1284,
   output        cfg_en1285,
   output        cfg_en1286,
   output        cfg_en1287,
   output        cfg_en1288,
   output        cfg_en1289,
   output        cfg_en1290,
   output        cfg_en1291,
   output        cfg_en1292,
   output        cfg_en1293,
   output        cfg_en1294,
   output        cfg_en1295,
   output        cfg_en1296,
   output        cfg_en1297,
   output        cfg_en1298,
   output        cfg_en1299,
   output        cfg_en1300,
   output        cfg_en1301,
   output        cfg_en1302,
   output        cfg_en1303,
   output        cfg_en1304,
   output        cfg_en1305,
   output        cfg_en1306,
   output        cfg_en1307,
   output        cfg_en1308,
   output        cfg_en1309,
   output        cfg_en1310,
   output        cfg_en1311,
   output        cfg_en1312,
   output        cfg_en1313,
   output        cfg_en1314,
   output        cfg_en1315,
   output        cfg_en1316,
   output        cfg_en1317,
   output        cfg_en1318,
   output        cfg_en1319,
   output        cfg_en1320,
   output        cfg_en1321,
   output        cfg_en1322,
   output        cfg_en1323,
   output        cfg_en1324,
   output        cfg_en1325,
   output        cfg_en1326,
   output        cfg_en1327,
   output        cfg_en1328,
   output        cfg_en1329,
   output        cfg_en1330,
   output        cfg_en1331,
   output        cfg_en1332,
   output        cfg_en1333,
   output        cfg_en1334,
   output        cfg_en1335,
   output        cfg_en1336,
   output        cfg_en1337,
   output        cfg_en1338,
   output        cfg_en1339,
   output        cfg_en1340,
   output        cfg_en1341,
   output        cfg_en1342,
   output        cfg_en1343,
   output        cfg_en1344,
   output        cfg_en1345,
   output        cfg_en1346,
   output        cfg_en1347,
   output        cfg_en1348,
   output        cfg_en1349,
   output        cfg_en1350,
   output        cfg_en1351,
   output        cfg_en1352,
   output        cfg_en1353,
   output        cfg_en1354,
   output        cfg_en1355,
   output        cfg_en1356,
   output        cfg_en1357,
   output        cfg_en1358,
   output        cfg_en1359,
   output        cfg_en1360,
   output        cfg_en1361,
   output        cfg_en1362,
   output        cfg_en1363,
   output        cfg_en1364,
   output        cfg_en1365,
   output        cfg_en1366,
   output        cfg_en1367,
   output        cfg_en1368,
   output        cfg_en1369,
   output        cfg_en1370,
   output        cfg_en1371,
   output        cfg_en1372,
   output        cfg_en1373,
   output        cfg_en1374,
   output        cfg_en1375,
   output        cfg_en1376,
   output        cfg_en1377,
   output        cfg_en1378,
   output        cfg_en1379,
   output        cfg_en1380,
   output        cfg_en1381,
   output        cfg_en1382,
   output        cfg_en1383,
   output        cfg_en1384,
   output        cfg_en1385,
   output        cfg_en1386,
   output        cfg_en1387,
   output        cfg_en1388,
   output        cfg_en1389,
   output        cfg_en1390,
   output        cfg_en1391,
   output        cfg_en1392,
   output        cfg_en1393,
   output        cfg_en1394,
   output        cfg_en1395,
   output        cfg_en1396,
   output        cfg_en1397,
   output        cfg_en1398,
   output        cfg_en1399,
   output        cfg_en1400,
   output        cfg_en1401,
   output        cfg_en1402,
   output        cfg_en1403,
   output        cfg_en1404,
   output        cfg_en1405,
   output        cfg_en1406,
   output        cfg_en1407,
   output        cfg_en1408,
   output        cfg_en1409,
   output        cfg_en1410,
   output        cfg_en1411,
   output        cfg_en1412,
   output        cfg_en1413,
   output        cfg_en1414,
   output        cfg_en1415,
   output        cfg_en1416,
   output        cfg_en1417,
   output        cfg_en1418,
   output        cfg_en1419,
   output        cfg_en1420,
   output        cfg_en1421,
   output        cfg_en1422,
   output        cfg_en1423,
   output        cfg_en1424,
   output        cfg_en1425,
   output        cfg_en1426,
   output        cfg_en1427,
   output        cfg_en1428,
   output        cfg_en1429,
   output        cfg_en1430,
   output        cfg_en1431,
   output        cfg_en1432,
   output        cfg_en1433,
   output        cfg_en1434,
   output        cfg_en1435,
   output        cfg_en1436,
   output        cfg_en1437,
   output        cfg_en1438,
   output        cfg_en1439,
   output        cfg_en1440,
   output        cfg_en1441,
   output        cfg_en1442,
   output        cfg_en1443,
   output        cfg_en1444,
   output        cfg_en1445,
   output        cfg_en1446,
   output        cfg_en1447,
   output        cfg_en1448,
   output        cfg_en1449,
   output        cfg_en1450,
   output        cfg_en1451,
   output        cfg_en1452,
   output        cfg_en1453,
   output        cfg_en1454,
   output        cfg_en1455,
   output        cfg_en1456,
   output        cfg_en1457,
   output        cfg_en1458,
   output        cfg_en1459,
   output        cfg_en1460,
   output        cfg_en1461,
   output        cfg_en1462,
   output        cfg_en1463,
   output        cfg_en1464,
   output        cfg_en1465,
   output        cfg_en1466,
   output        cfg_en1467,
   output        cfg_en1468,
   output        cfg_en1469,
   output        cfg_en1470,
   output        cfg_en1471,
   output        cfg_en1472,
   output        cfg_en1473,
   output        cfg_en1474,
   output        cfg_en1475,
   output        cfg_en1476,
   output        cfg_en1477,
   output        cfg_en1478,
   output        cfg_en1479,
   output        cfg_en1480,
   output        cfg_en1481,
   output        cfg_en1482,
   output        cfg_en1483,
   output        cfg_en1484,
   output        cfg_en1485,
   output        cfg_en1486,
   output        cfg_en1487,
   output        cfg_en1488,
   output        cfg_en1489,
   output        cfg_en1490,
   output        cfg_en1491,
   output        cfg_en1492,
   output        cfg_en1493,
   output        cfg_en1494,
   output        cfg_en1495,
   output        cfg_en1496,
   output        cfg_en1497,
   output        cfg_en1498,
   output        cfg_en1499,
   output        cfg_en1500,
   output        cfg_en1501,
   output        cfg_en1502,
   output        cfg_en1503,
   output        cfg_en1504,
   output        cfg_en1505,
   output        cfg_en1506,
   output        cfg_en1507,
   output        cfg_en1508,
   output        cfg_en1509,
   output        cfg_en1510,
   output        cfg_en1511,
   output        cfg_en1512,
   output        cfg_en1513,
   output        cfg_en1514,
   output        cfg_en1515,
   output        cfg_en1516,
   output        cfg_en1517,
   output        cfg_en1518,
   output        cfg_en1519,
   output        cfg_en1520,
   output        cfg_en1521,
   output        cfg_en1522,
   output        cfg_en1523,
   output        cfg_en1524,
   output        cfg_en1525,
   output        cfg_en1526,
   output        cfg_en1527,
   output        cfg_en1528,
   output        cfg_en1529,
   output        cfg_en1530,
   output        cfg_en1531,
   output        cfg_en1532,
   output        cfg_en1533,
   output        cfg_en1534,
   output        cfg_en1535,
   output        cfg_en1536,
   output        cfg_en1537,
   output        cfg_en1538,
   output        cfg_en1539,
   output        cfg_en1540,
   output        cfg_en1541,
   output        cfg_en1542,
   output        cfg_en1543,
   output        cfg_en1544,
   output        cfg_en1545,
   output        cfg_en1546,
   output        cfg_en1547,
   output        cfg_en1548,
   output        cfg_en1549,
   output        cfg_en1550,
   output        cfg_en1551,
   output        cfg_en1552,
   output        cfg_en1553,
   output        cfg_en1554,
   output        cfg_en1555,
   output        cfg_en1556,
   output        cfg_en1557,
   output        cfg_en1558,
   output        cfg_en1559,
   output        cfg_en1560,
   output        cfg_en1561,
   output        cfg_en1562,
   output        cfg_en1563,
   output        cfg_en1564,
   output        cfg_en1565,
   output        cfg_en1566,
   output        cfg_en1567,
   output        cfg_en1568,
   output        cfg_en1569,
   output        cfg_en1570,
   output        cfg_en1571,
   output        cfg_en1572,
   output        cfg_en1573,
   output        cfg_en1574,
   output        cfg_en1575,
   output        cfg_en1576,
   output        cfg_en1577,
   output        cfg_en1578,
   output        cfg_en1579,
   output        cfg_en1580,
   output        cfg_en1581,
   output        cfg_en1582,
   output        cfg_en1583,
   output        cfg_en1584,
   output        cfg_en1585,
   output        cfg_en1586,
   output        cfg_en1587,
   output        cfg_en1588,
   output        cfg_en1589,
   output        cfg_en1590,
   output        cfg_en1591,
   output        cfg_en1592,
   output        cfg_en1593,
   output        cfg_en1594,
   output        cfg_en1595,
   output        cfg_en1596,
   output        cfg_en1597,
   output        cfg_en1598,
   output        cfg_en1599,
   output        cfg_en1600,
   output        cfg_en1601,
   output        cfg_en1602,
   output        cfg_en1603,
   output        cfg_en1604,
   output        cfg_en1605,
   output        cfg_en1606,
   output        cfg_en1607,
   output        cfg_en1608,
   output        cfg_en1609,
   output        cfg_en1610,
   output        cfg_en1611,
   output        cfg_en1612,
   output        cfg_en1613,
   output        cfg_en1614,
   output        cfg_en1615,
   output        cfg_en1616,
   output        cfg_en1617,
   output        cfg_en1618,
   output        cfg_en1619,
   output        cfg_en1620,
   output        cfg_en1621,
   output        cfg_en1622,
   output        cfg_en1623,
   output        cfg_en1624,
   output        cfg_en1625,
   output        cfg_en1626,
   output        cfg_en1627,
   output        cfg_en1628,
   output        cfg_en1629,
   output        cfg_en1630,
   output        cfg_en1631,
   output        cfg_en1632,
   output        cfg_en1633,
   output        cfg_en1634,
   output        cfg_en1635,
   output        cfg_en1636,
   output        cfg_en1637,
   output        cfg_en1638,
   output        cfg_en1639,
   output        cfg_en1640,
   output        cfg_en1641,
   output        cfg_en1642,
   output        cfg_en1643,
   output        cfg_en1644,
   output        cfg_en1645,
   output        cfg_en1646,
   output        cfg_en1647,
   output        cfg_en1648,
   output        cfg_en1649,
   output        cfg_en1650,
   output        cfg_en1651,
   output        cfg_en1652,
   output        cfg_en1653,
   output        cfg_en1654,
   output        cfg_en1655,
   output        cfg_en1656,
   output        cfg_en1657,
   output        cfg_en1658,
   output        cfg_en1659,
   output        cfg_en1660,
   output        cfg_en1661,
   output        cfg_en1662,
   output        cfg_en1663,
   output        cfg_en1664,
   output        cfg_en1665,
   output        cfg_en1666,
   output        cfg_en1667,
   output        cfg_en1668,
   output        cfg_en1669,
   output        cfg_en1670,
   output        cfg_en1671,
   output        cfg_en1672,
   output        cfg_en1673,
   output        cfg_en1674,
   output        cfg_en1675,
   output        cfg_en1676,
   output        cfg_en1677,
   output        cfg_en1678,
   output        cfg_en1679,
   output        cfg_en1680,
   output        cfg_en1681,
   output        cfg_en1682,
   output        cfg_en1683,
   output        cfg_en1684,
   output        cfg_en1685,
   output        cfg_en1686,
   output        cfg_en1687,
   output        cfg_en1688,
   output        cfg_en1689,
   output        cfg_en1690,
   output        cfg_en1691,
   output        cfg_en1692,
   output        cfg_en1693,
   output        cfg_en1694,
   output        cfg_en1695,
   output        cfg_en1696,
   output        cfg_en1697,
   output        cfg_en1698,
   output        cfg_en1699,
   output        cfg_en1700,
   output        cfg_en1701,
   output        cfg_en1702,
   output        cfg_en1703,
   output        cfg_en1704,
   output        cfg_en1705,
   output        cfg_en1706,
   output        cfg_en1707,
   output        cfg_en1708,
   output        cfg_en1709,
   output        cfg_en1710,
   output        cfg_en1711,
   output        cfg_en1712,
   output        cfg_en1713,
   output        cfg_en1714,
   output        cfg_en1715,
   output        cfg_en1716,
   output        cfg_en1717,
   output        cfg_en1718,
   output        cfg_en1719,
   output        cfg_en1720,
   output        cfg_en1721,
   output        cfg_en1722,
   output        cfg_en1723,
   output        cfg_en1724,
   output        cfg_en1725,
   output        cfg_en1726,
   output        cfg_en1727,
   output        cfg_en1728,
   output        cfg_en1729,
   output        cfg_en1730,
   output        cfg_en1731,
   output        cfg_en1732,
   output        cfg_en1733,
   output        cfg_en1734,
   output        cfg_en1735,
   output        cfg_en1736,
   output        cfg_en1737,
   output        cfg_en1738,
   output        cfg_en1739,
   output        cfg_en1740,
   output        cfg_en1741,
   output        cfg_en1742,
   output        cfg_en1743,
   output        cfg_en1744,
   output        cfg_en1745,
   output        cfg_en1746,
   output        cfg_en1747,
   output        cfg_en1748,
   output        cfg_en1749,
   output        cfg_en1750,
   output        cfg_en1751,
   output        cfg_en1752,
   output        cfg_en1753,
   output        cfg_en1754,
   output        cfg_en1755,
   output        cfg_en1756,
   output        cfg_en1757,
   output        cfg_en1758,
   output        cfg_en1759,
   output        cfg_en1760,
   output        cfg_en1761,
   output        cfg_en1762,
   output        cfg_en1763,
   output        cfg_en1764,
   output        cfg_en1765,
   output        cfg_en1766,
   output        cfg_en1767,
   output        cfg_en1768,
   output        cfg_en1769,
   output        cfg_en1770,
   output        cfg_en1771,
   output        cfg_en1772,
   output        cfg_en1773,
   output        cfg_en1774,
   output        cfg_en1775,
   output        cfg_en1776,
   output        cfg_en1777,
   output        cfg_en1778,
   output        cfg_en1779,
   output        cfg_en1780,
   output        cfg_en1781,
   output        cfg_en1782,
   output        cfg_en1783,
   output        cfg_en1784,
   output        cfg_en1785,
   output        cfg_en1786,
   output        cfg_en1787,
   output        cfg_en1788,
   output        cfg_en1789,
   output        cfg_en1790,
   output        cfg_en1791,
   output        cfg_en1792,
   output        cfg_en1793,
   output        cfg_en1794,
   output        cfg_en1795,
   output        cfg_en1796,
   output        cfg_en1797,
   output        cfg_en1798,
   output        cfg_en1799,
   output        cfg_en1800,
   output        cfg_en1801,
   output        cfg_en1802,
   output        cfg_en1803,
   output        cfg_en1804,
   output        cfg_en1805,
   output        cfg_en1806,
   output        cfg_en1807,
   output        cfg_en1808,
   output        cfg_en1809,
   output        cfg_en1810,
   output        cfg_en1811,
   output        cfg_en1812,
   output        cfg_en1813,
   output        cfg_en1814,
   output        cfg_en1815,
   output        cfg_en1816,
   output        cfg_en1817,
   output        cfg_en1818,
   output        cfg_en1819,
   output        cfg_en1820,
   output        cfg_en1821,
   output        cfg_en1822,
   output        cfg_en1823,
   output        cfg_en1824,
   output        cfg_en1825,
   output        cfg_en1826,
   output        cfg_en1827,
   output        cfg_en1828,
   output        cfg_en1829,
   output        cfg_en1830,
   output        cfg_en1831,
   output        cfg_en1832,
   output        cfg_en1833,
   output        cfg_en1834,
   output        cfg_en1835,
   output        cfg_en1836,
   output        cfg_en1837,
   output        cfg_en1838,
   output        cfg_en1839,
   output        cfg_en1840,
   output        cfg_en1841,
   output        cfg_en1842,
   output        cfg_en1843,
   output        cfg_en1844,
   output        cfg_en1845,
   output        cfg_en1846,
   output        cfg_en1847,
   output        cfg_en1848,
   output        cfg_en1849,
   output        cfg_en1850,
   output        cfg_en1851,
   output        cfg_en1852,
   output        cfg_en1853,
   output        cfg_en1854,
   output        cfg_en1855,
   output        cfg_en1856,
   output        cfg_en1857,
   output        cfg_en1858,
   output        cfg_en1859,
   output        cfg_en1860,
   output        cfg_en1861,
   output        cfg_en1862,
   output        cfg_en1863,
   output        cfg_en1864,
   output        cfg_en1865,
   output        cfg_en1866,
   output        cfg_en1867,
   output        cfg_en1868,
   output        cfg_en1869,
   output        cfg_en1870,
   output        cfg_en1871,
   output        cfg_en1872,
   output        cfg_en1873,
   output        cfg_en1874,
   output        cfg_en1875,
   output        cfg_en1876,
   output        cfg_en1877,
   output        cfg_en1878,
   output        cfg_en1879,
   output        cfg_en1880,
   output        cfg_en1881,
   output        cfg_en1882,
   output        cfg_en1883,
   output        cfg_en1884,
   output        cfg_en1885,
   output        cfg_en1886,
   output        cfg_en1887,
   output        cfg_en1888,
   output        cfg_en1889,
   output        cfg_en1890,
   output        cfg_en1891,
   output        cfg_en1892,
   output        cfg_en1893,
   output        cfg_en1894,
   output        cfg_en1895,
   output        cfg_en1896,
   output        cfg_en1897,
   output        cfg_en1898,
   output        cfg_en1899,
   output        cfg_en1900,
   output        cfg_en1901,
   output        cfg_en1902,
   output        cfg_en1903,
   output        cfg_en1904,
   output        cfg_en1905,
   output        cfg_en1906,
   output        cfg_en1907,
   output        cfg_en1908,
   output        cfg_en1909,
   output        cfg_en1910,
   output        cfg_en1911,
   output        cfg_en1912,
   output        cfg_en1913,
   output        cfg_en1914,
   output        cfg_en1915,
   output        cfg_en1916,
   output        cfg_en1917,
   output        cfg_en1918,
   output        cfg_en1919,
   output        cfg_en1920,
   output        cfg_en1921,
   output        cfg_en1922,
   output        cfg_en1923,
   output        cfg_en1924,
   output        cfg_en1925,
   output        cfg_en1926,
   output        cfg_en1927,
   output        cfg_en1928,
   output        cfg_en1929,
   output        cfg_en1930,
   output        cfg_en1931,
   output        cfg_en1932,
   output        cfg_en1933,
   output        cfg_en1934,
   output        cfg_en1935,
   output        cfg_en1936,
   output        cfg_en1937,
   output        cfg_en1938,
   output        cfg_en1939,
   output        cfg_en1940,
   output        cfg_en1941,
   output        cfg_en1942,
   output        cfg_en1943,
   output        cfg_en1944,
   output        cfg_en1945,
   output        cfg_en1946,
   output        cfg_en1947,
   output        cfg_en1948,
   output        cfg_en1949,
   output        cfg_en1950,
   output        cfg_en1951,
   output        cfg_en1952,
   output        cfg_en1953,
   output        cfg_en1954,
   output        cfg_en1955,
   output        cfg_en1956,
   output        cfg_en1957,
   output        cfg_en1958,
   output        cfg_en1959,
   output        cfg_en1960,
   output        cfg_en1961,
   output        cfg_en1962,
   output        cfg_en1963,
   output        cfg_en1964,
   output        cfg_en1965,
   output        cfg_en1966,
   output        cfg_en1967,
   output        cfg_en1968,
   output        cfg_en1969,
   output        cfg_en1970,
   output        cfg_en1971,
   output        cfg_en1972,
   output        cfg_en1973,
   output        cfg_en1974,
   output        cfg_en1975,
   output        cfg_en1976,
   output        cfg_en1977,
   output        cfg_en1978,
   output        cfg_en1979,
   output        cfg_en1980,
   output        cfg_en1981,
   output        cfg_en1982,
   output        cfg_en1983,
   output        cfg_en1984,
   output        cfg_en1985,
   output        cfg_en1986,
   output        cfg_en1987,
   output        cfg_en1988,
   output        cfg_en1989,
   output        cfg_en1990,
   output        cfg_en1991,
   output        cfg_en1992,
   output        cfg_en1993,
   output        cfg_en1994,
   output        cfg_en1995,
   output        cfg_en1996,
   output        cfg_en1997,
   output        cfg_en1998,
   output        cfg_en1999,
   output        cfg_en2000,
   output        cfg_en2001,
   output        cfg_en2002,
   output        cfg_en2003,
   output        cfg_en2004,
   output        cfg_en2005,
   output        cfg_en2006,
   output        cfg_en2007,
   output        cfg_en2008,
   output        cfg_en2009,
   output        cfg_en2010,
   output        cfg_en2011,
   output        cfg_en2012,
   output        cfg_en2013,
   output        cfg_en2014,
   output        cfg_en2015,
   output        cfg_en2016,
   output        cfg_en2017,
   output        cfg_en2018,
   output        cfg_en2019,
   output        cfg_en2020,
   output        cfg_en2021,
   output        cfg_en2022,
   output        cfg_en2023,
   output        cfg_en2024,
   output        cfg_en2025,
   output        cfg_en2026,
   output        cfg_en2027,
   output        cfg_en2028,
   output        cfg_en2029,
   output        cfg_en2030,
   output        cfg_en2031,
   output        cfg_en2032,
   output        cfg_en2033,
   output        cfg_en2034,
   output        cfg_en2035,
   output        cfg_en2036,
   output        cfg_en2037,
   output        cfg_en2038,
   output        cfg_en2039,
   output        cfg_en2040,
   output        cfg_en2041,
   output        cfg_en2042,
   output        cfg_en2043,
   output        cfg_en2044,
   output        cfg_en2045,
   output        cfg_en2046,
   output        cfg_en2047,
   output        cfg_en2048,
   output        cfg_en2049,
   output        cfg_en2050,
   output        cfg_en2051,
   output        cfg_en2052,
   output        cfg_en2053,
   output        cfg_en2054,
   output        cfg_en2055,
   output        cfg_en2056,
   output        cfg_en2057,
   output        cfg_en2058,
   output        cfg_en2059,
   output        cfg_en2060,
   output        cfg_en2061,
   output        cfg_en2062,
   output        cfg_en2063,
   output        cfg_en2064,
   output        cfg_en2065,
   output        cfg_en2066,
   output        cfg_en2067,
   output        cfg_en2068,
   output        cfg_en2069,
   output        cfg_en2070,
   output        cfg_en2071,
   output        cfg_en2072,
   output        cfg_en2073,
   output        cfg_en2074,
   output        cfg_en2075,
   output        cfg_en2076,
   output        cfg_en2077,
   output        cfg_en2078,
   output        cfg_en2079,
   output        cfg_en2080,
   output        cfg_en2081,
   output        cfg_en2082,
   output        cfg_en2083,
   output        cfg_en2084,
   output        cfg_en2085,
   output        cfg_en2086,
   output        cfg_en2087,
   output        cfg_en2088,
   output        cfg_en2089,
   output        cfg_en2090,
   output        cfg_en2091,
   output        cfg_en2092,
   output        cfg_en2093,
   output        cfg_en2094,
   output        cfg_en2095,
   output        cfg_en2096,
   output        cfg_en2097,
   output        cfg_en2098,
   output        cfg_en2099,
   output        cfg_en2100,
   output        cfg_en2101,
   output        cfg_en2102,
   output        cfg_en2103,
   output        cfg_en2104,
   output        cfg_en2105,
   output        cfg_en2106,
   output        cfg_en2107,
   output        cfg_en2108,
   output        cfg_en2109,
   output        cfg_en2110,
   output        cfg_en2111,
   output        cfg_en2112,
   output        cfg_en2113,
   output        cfg_en2114,
   output        cfg_en2115,
   output        cfg_en2116,
   output        cfg_en2117,
   output        cfg_en2118,
   output        cfg_en2119,
   output        cfg_en2120,
   output        cfg_en2121,
   output        cfg_en2122,
   output        cfg_en2123,
   output        cfg_en2124,
   output        cfg_en2125,
   output        cfg_en2126,
   output        cfg_en2127,
   output        cfg_en2128,
   output        cfg_en2129,
   output        cfg_en2130,
   output        cfg_en2131,
   output        cfg_en2132,
   output        cfg_en2133,
   output        cfg_en2134,
   output        cfg_en2135,
   output        cfg_en2136,
   output        cfg_en2137,
   output        cfg_en2138,
   output        cfg_en2139,
   output        cfg_en2140,
   output        cfg_en2141,
   output        cfg_en2142,
   output        cfg_en2143,
   output        cfg_en2144,
   output        cfg_en2145,
   output        cfg_en2146,
   output        cfg_en2147,
   output        cfg_en2148,
   output        cfg_en2149,
   output        cfg_en2150,
   output        cfg_en2151,
   output        cfg_en2152,
   output        cfg_en2153,
   output        cfg_en2154,
   output        cfg_en2155,
   output        cfg_en2156,
   output        cfg_en2157,
   output        cfg_en2158,
   output        cfg_en2159,
   output        cfg_en2160,
   output        cfg_en2161,
   output        cfg_en2162,
   output        cfg_en2163,
   output        cfg_en2164,
   output        cfg_en2165,
   output        cfg_en2166,
   output        cfg_en2167,
   output        cfg_en2168,
   output        cfg_en2169,
   output        cfg_en2170,
   output        cfg_en2171,
   output        cfg_en2172,
   output        cfg_en2173,
   output        cfg_en2174,
   output        cfg_en2175,
   output        cfg_en2176,
   output        cfg_en2177,
   output        cfg_en2178,
   output        cfg_en2179,
   output        cfg_en2180,
   output        cfg_en2181,
   output        cfg_en2182,
   output        cfg_en2183,
   output        cfg_en2184,
   output        cfg_en2185,
   output        cfg_en2186,
   output        cfg_en2187,
   output        cfg_en2188,
   output        cfg_en2189,
   output        cfg_en2190,
   output        cfg_en2191,
   output        cfg_en2192,
   output        cfg_en2193,
   output        cfg_en2194,
   output        cfg_en2195,
   output        cfg_en2196,
   output        cfg_en2197,
   output        cfg_en2198,
   output        cfg_en2199,
   output        cfg_en2200,
   output        cfg_en2201,
   output        cfg_en2202,
   output        cfg_en2203,
   output        cfg_en2204,
   output        cfg_en2205,
   output        cfg_en2206,
   output        cfg_en2207,
   output        cfg_en2208,
   output        cfg_en2209,
   output        cfg_en2210,
   output        cfg_en2211,
   output        cfg_en2212,
   output        cfg_en2213,
   output        cfg_en2214,
   output        cfg_en2215,
   output        cfg_en2216,
   output        cfg_en2217,
   output        cfg_en2218,
   output        cfg_en2219,
   output        cfg_en2220,
   output        cfg_en2221,
   output        cfg_en2222,
   output        cfg_en2223,
   output        cfg_en2224,
   output        cfg_en2225,
   output        cfg_en2226,
   output        cfg_en2227,
   output        cfg_en2228,
   output        cfg_en2229,
   output        cfg_en2230,
   output        cfg_en2231,
   output        cfg_en2232,
   output        cfg_en2233,
   output        cfg_en2234,
   output        cfg_en2235,
   output        cfg_en2236,
   output        cfg_en2237,
   output        cfg_en2238,
   output        cfg_en2239,
   output        cfg_en2240,
   output        cfg_en2241,
   output        cfg_en2242,
   output        cfg_en2243,
   output        cfg_en2244,
   output        cfg_en2245,
   output        cfg_en2246,
   output        cfg_en2247,
   output        cfg_en2248,
   output        cfg_en2249,
   output        cfg_en2250,
   output        cfg_en2251,
   output        cfg_en2252,
   output        cfg_en2253,
   output        cfg_en2254,
   output        cfg_en2255,
   output        cfg_en2256,
   output        cfg_en2257,
   output        cfg_en2258,
   output        cfg_en2259,
   output        cfg_en2260,
   output        cfg_en2261,
   output        cfg_en2262,
   output        cfg_en2263,
   output        cfg_en2264,
   output        cfg_en2265,
   output        cfg_en2266,
   output        cfg_en2267,
   output        cfg_en2268,
   output        cfg_en2269,
   output        cfg_en2270,
   output        cfg_en2271,
   output        cfg_en2272,
   output        cfg_en2273,
   output        cfg_en2274,
   output        cfg_en2275,
   output        cfg_en2276,
   output        cfg_en2277,
   output        cfg_en2278,
   output        cfg_en2279,
   output        cfg_en2280,
   output        cfg_en2281,
   output        cfg_en2282,
   output        cfg_en2283,
   output        cfg_en2284,
   output        cfg_en2285,
   output        cfg_en2286,
   output        cfg_en2287,
   output        cfg_en2288,
   output        cfg_en2289,
   output        cfg_en2290,
   output        cfg_en2291,
   output        cfg_en2292,
   output        cfg_en2293,
   output        cfg_en2294,
   output        cfg_en2295,
   output        cfg_en2296,
   output        cfg_en2297,
   output        cfg_en2298,
   output        cfg_en2299,
   output        cfg_en2300,
   output        cfg_en2301,
   output        cfg_en2302,
   output        cfg_en2303,
   output        cfg_en2304,
   output        cfg_en2305,
   output        cfg_en2306,
   output        cfg_en2307,
   output        cfg_en2308,
   output        cfg_en2309,
   output        cfg_en2310,
   output        cfg_en2311,
   output        cfg_en2312,
   output        cfg_en2313,
   output        cfg_en2314,
   output        cfg_en2315,
   output        cfg_en2316,
   output        cfg_en2317,
   output        cfg_en2318,
   output        cfg_en2319,
   output        cfg_en2320,
   output        cfg_en2321,
   output        cfg_en2322,
   output        cfg_en2323,
   output        cfg_en2324,
   output        cfg_en2325,
   output        cfg_en2326,
   output        cfg_en2327,
   output        cfg_en2328,
   output        cfg_en2329,
   output        cfg_en2330,
   output        cfg_en2331,
   output        cfg_en2332,
   output        cfg_en2333,
   output        cfg_en2334,
   output        cfg_en2335,
   output        cfg_en2336,
   output        cfg_en2337,
   output        cfg_en2338,
   output        cfg_en2339,
   output        cfg_en2340,
   output        cfg_en2341,
   output        cfg_en2342,
   output        cfg_en2343,
   output        cfg_en2344,
   output        cfg_en2345,
   output        cfg_en2346,
   output        cfg_en2347,
   output        cfg_en2348,
   output        cfg_en2349,
   output        cfg_en2350,
   output        cfg_en2351,
   output        cfg_en2352,
   output        cfg_en2353,
   output        cfg_en2354,
   output        cfg_en2355,
   output        cfg_en2356,
   output        cfg_en2357,
   output        cfg_en2358,
   output        cfg_en2359,
   output        cfg_en2360,
   output        cfg_en2361,
   output        cfg_en2362,
   output        cfg_en2363,
   output        cfg_en2364,
   output        cfg_en2365,
   output        cfg_en2366,
   output        cfg_en2367,
   output        cfg_en2368,
   output        cfg_en2369,
   output        cfg_en2370,
   output        cfg_en2371,
   output        cfg_en2372,
   output        cfg_en2373,
   output        cfg_en2374,
   output        cfg_en2375,
   output        cfg_en2376,
   output        cfg_en2377,
   output        cfg_en2378,
   output        cfg_en2379,
   output        cfg_en2380,
   output        cfg_en2381,
   output        cfg_en2382,
   output        cfg_en2383,
   output        cfg_en2384,
   output        cfg_en2385,
   output        cfg_en2386,
   output        cfg_en2387,
   output        cfg_en2388,
   output        cfg_en2389,
   output        cfg_en2390,
   output        cfg_en2391,
   output        cfg_en2392,
   output        cfg_en2393,
   output        cfg_en2394,
   output        cfg_en2395,
   output        cfg_en2396,
   output        cfg_en2397,
   output        cfg_en2398,
   output        cfg_en2399,
   output        cfg_en2400,
   output        cfg_en2401,
   output        cfg_en2402,
   output        cfg_en2403,
   output        cfg_en2404,
   output        cfg_en2405,
   output        cfg_en2406,
   output        cfg_en2407,
   output        cfg_en2408,
   output        cfg_en2409,
   output        cfg_en2410,
   output        cfg_en2411,
   output        cfg_en2412,
   output        cfg_en2413,
   output        cfg_en2414,
   output        cfg_en2415,
   output        cfg_en2416,
   output        cfg_en2417,
   output        cfg_en2418,
   output        cfg_en2419,
   output        cfg_en2420,
   output        cfg_en2421,
   output        cfg_en2422,
   output        cfg_en2423,
   output        cfg_en2424,
   output        cfg_en2425,
   output        cfg_en2426,
   output        cfg_en2427,
   output        cfg_en2428,
   output        cfg_en2429,
   output        cfg_en2430,
   output        cfg_en2431,
   output        cfg_en2432,
   output        cfg_en2433,
   output        cfg_en2434,
   output        cfg_en2435,
   output        cfg_en2436,
   output        cfg_en2437,
   output        cfg_en2438,
   output        cfg_en2439,
   output        cfg_en2440,
   output        cfg_en2441,
   output        cfg_en2442,
   output        cfg_en2443,
   output        cfg_en2444,
   output        cfg_en2445,
   output        cfg_en2446,
   output        cfg_en2447,
   output        cfg_en2448,
   output        cfg_en2449,
   output        cfg_en2450,
   output        cfg_en2451,
   output        cfg_en2452,
   output        cfg_en2453,
   output        cfg_en2454,
   output        cfg_en2455,
   output        cfg_en2456,
   output        cfg_en2457,
   output        cfg_en2458,
   output        cfg_en2459,
   output        cfg_en2460,
   output        cfg_en2461,
   output        cfg_en2462,
   output        cfg_en2463,
   output        cfg_en2464,
   output        cfg_en2465,
   output        cfg_en2466,
   output        cfg_en2467,
   output        cfg_en2468,
   output        cfg_en2469,
   output        cfg_en2470,
   output        cfg_en2471,
   output        cfg_en2472,
   output        cfg_en2473,
   output        cfg_en2474,
   output        cfg_en2475,
   output        cfg_en2476,
   output        cfg_en2477,
   output        cfg_en2478,
   output        cfg_en2479,
   output        cfg_en2480,
   output        cfg_en2481,
   output        cfg_en2482,
   output        cfg_en2483,
   output        cfg_en2484,
   output        cfg_en2485,
   output        cfg_en2486,
   output        cfg_en2487,
   output        cfg_en2488,
   output        cfg_en2489,
   output        cfg_en2490,
   output        cfg_en2491,
   output        cfg_en2492,
   output        cfg_en2493,
   output        cfg_en2494,
   output        cfg_en2495,
   output        cfg_en2496,
   output        cfg_en2497,
   output        cfg_en2498,
   output        cfg_en2499,
   output        cfg_en2500,
   output        cfg_en2501,
   output        cfg_en2502,
   output        cfg_en2503,
   output        cfg_en2504,
   output        cfg_en2505,
   output        cfg_en2506,
   output        cfg_en2507,
   output        cfg_en2508,
   output        cfg_en2509,
   output        cfg_en2510,
   output        cfg_en2511,
   output        cfg_en2512,
   output        cfg_en2513,
   output        cfg_en2514,
   output        cfg_en2515,
   output        cfg_en2516,
   output        cfg_en2517,
   output        cfg_en2518,
   output        cfg_en2519,
   output        cfg_en2520,
   output        cfg_en2521,
   output        cfg_en2522,
   output        cfg_en2523,
   output        cfg_en2524,
   output        cfg_en2525,
   output        cfg_en2526,
   output        cfg_en2527,
   output        cfg_en2528,
   output        cfg_en2529,
   output        cfg_en2530,
   output        cfg_en2531,
   output        cfg_en2532,
   output        cfg_en2533,
   output        cfg_en2534,
   output        cfg_en2535,
   output        cfg_en2536,
   output        cfg_en2537,
   output        cfg_en2538,
   output        cfg_en2539,
   output        cfg_en2540,
   output        cfg_en2541,
   output        cfg_en2542,
   output        cfg_en2543,
   output        cfg_en2544,
   output        cfg_en2545,
   output        cfg_en2546,
   output        cfg_en2547,
   output        cfg_en2548,
   output        cfg_en2549,
   output        cfg_en2550,
   output        cfg_en2551,
   output        cfg_en2552,
   output        cfg_en2553,
   output        cfg_en2554,
   output        cfg_en2555,
   output        cfg_en2556,
   output        cfg_en2557,
   output        cfg_en2558,
   output        cfg_en2559,
   output        cfg_en2560,
   output        cfg_en2561,
   output        cfg_en2562,
   output        cfg_en2563,
   output        cfg_en2564,
   output        cfg_en2565,
   output        cfg_en2566,
   output        cfg_en2567,
   output        cfg_en2568,
   output        cfg_en2569,
   output        cfg_en2570,
   output        cfg_en2571,
   output        cfg_en2572,
   output        cfg_en2573,
   output        cfg_en2574,
   output        cfg_en2575,
   output        cfg_en2576,
   output        cfg_en2577,
   output        cfg_en2578,
   output        cfg_en2579,
   output        cfg_en2580,
   output        cfg_en2581,
   output        cfg_en2582,
   output        cfg_en2583,
   output        cfg_en2584,
   output        cfg_en2585,
   output        cfg_en2586,
   output        cfg_en2587,
   output        cfg_en2588,
   output        cfg_en2589,
   output        cfg_en2590,
   output        cfg_en2591,
   output        cfg_en2592,
   output        cfg_en2593,
   output        cfg_en2594,
   output        cfg_en2595,
   output        cfg_en2596,
   output        cfg_en2597,
   output        cfg_en2598,
   output        cfg_en2599,
   output        cfg_en2600,
   output        cfg_en2601,
   output        cfg_en2602,
   output        cfg_en2603,
   output        cfg_en2604,
   output        cfg_en2605,
   output        cfg_en2606,
   output        cfg_en2607,
   output        cfg_en2608,
   output        cfg_en2609,
   output        cfg_en2610,
   output        cfg_en2611,
   output        cfg_en2612,
   output        cfg_en2613,
   output        cfg_en2614,
   output        cfg_en2615,
   output        cfg_en2616,
   output        cfg_en2617,
   output        cfg_en2618,
   output        cfg_en2619,
   output        cfg_en2620,
   output        cfg_en2621,
   output        cfg_en2622,
   output        cfg_en2623,
   output        cfg_en2624,
   output        cfg_en2625,
   output        cfg_en2626,
   output        cfg_en2627,
   output        cfg_en2628,
   output        cfg_en2629,
   output        cfg_en2630,
   output        cfg_en2631,
   output        cfg_en2632,
   output        cfg_en2633,
   output        cfg_en2634,
   output        cfg_en2635,
   output        cfg_en2636,
   output        cfg_en2637,
   output        cfg_en2638,
   output        cfg_en2639,
   output        cfg_en2640,
   output        cfg_en2641,
   output        cfg_en2642,
   output        cfg_en2643,
   output        cfg_en2644,
   output        cfg_en2645,
   output        cfg_en2646,
   output        cfg_en2647,
   output        cfg_en2648,
   output        cfg_en2649,
   output        cfg_en2650,
   output        cfg_en2651,
   output        cfg_en2652,
   output        cfg_en2653,
   output        cfg_en2654,
   output        cfg_en2655,
   output        cfg_en2656,
   output        cfg_en2657,
   output        cfg_en2658,
   output        cfg_en2659,
   output        cfg_en2660,
   output        cfg_en2661,
   output        cfg_en2662,
   output        cfg_en2663,
   output        cfg_en2664,
   output        cfg_en2665,
   output        cfg_en2666,
   output        cfg_en2667,
   output        cfg_en2668,
   output        cfg_en2669,
   output        cfg_en2670,
   output        cfg_en2671,
   output        cfg_en2672,
   output        cfg_en2673,
   output        cfg_en2674,
   output        cfg_en2675,
   output        cfg_en2676,
   output        cfg_en2677,
   output        cfg_en2678,
   output        cfg_en2679,
   output        cfg_en2680,
   output        cfg_en2681,
   output        cfg_en2682,
   output        cfg_en2683,
   output        cfg_en2684,
   output        cfg_en2685,
   output        cfg_en2686,
   output        cfg_en2687,
   output        cfg_en2688,
   output        cfg_en2689,
   output        cfg_en2690,
   output        cfg_en2691,
   output        cfg_en2692,
   output        cfg_en2693,
   output        cfg_en2694,
   output        cfg_en2695,
   output        cfg_en2696,
   output        cfg_en2697,
   output        cfg_en2698,
   output        cfg_en2699,
   output        cfg_en2700,
   output        cfg_en2701,
   output        cfg_en2702,
   output        cfg_en2703,
   output        cfg_en2704,
   output        cfg_en2705,
   output        cfg_en2706,
   output        cfg_en2707,
   output        cfg_en2708,
   output        cfg_en2709,
   output        cfg_en2710,
   output        cfg_en2711,
   output        cfg_en2712,
   output        cfg_en2713,
   output        cfg_en2714,
   output        cfg_en2715,
   output        cfg_en2716,
   output        cfg_en2717,
   output        cfg_en2718,
   output        cfg_en2719,
   output        cfg_en2720,
   output        cfg_en2721,
   output        cfg_en2722,
   output        cfg_en2723,
   output        cfg_en2724,
   output        cfg_en2725,
   output        cfg_en2726,
   output        cfg_en2727,
   output        cfg_en2728,
   output        cfg_en2729,
   output        cfg_en2730,
   output        cfg_en2731,
   output        cfg_en2732,
   output        cfg_en2733,
   output        cfg_en2734,
   output        cfg_en2735,
   output        cfg_en2736,
   output        cfg_en2737,
   output        cfg_en2738,
   output        cfg_en2739,
   output        cfg_en2740,
   output        cfg_en2741,
   output        cfg_en2742,
   output        cfg_en2743,
   output        cfg_en2744,
   output        cfg_en2745,
   output        cfg_en2746,
   output        cfg_en2747,
   output        cfg_en2748,
   output        cfg_en2749,
   output        cfg_en2750,
   output        cfg_en2751,
   output        cfg_en2752,
   output        cfg_en2753,
   output        cfg_en2754,
   output        cfg_en2755,
   output        cfg_en2756,
   output        cfg_en2757,
   output        cfg_en2758,
   output        cfg_en2759,
   output        cfg_en2760,
   output        cfg_en2761,
   output        cfg_en2762,
   output        cfg_en2763,
   output        cfg_en2764,
   output        cfg_en2765,
   output        cfg_en2766,
   output        cfg_en2767,
   output        cfg_en2768,
   output        cfg_en2769,
   output        cfg_en2770,
   output        cfg_en2771,
   output        cfg_en2772,
   output        cfg_en2773,
   output        cfg_en2774,
   output        cfg_en2775,
   output        cfg_en2776,
   output        cfg_en2777,
   output        cfg_en2778,
   output        cfg_en2779,
   output        cfg_en2780,
   output        cfg_en2781,
   output        cfg_en2782,
   output        cfg_en2783,
   output        cfg_en2784,
   output        cfg_en2785,
   output        cfg_en2786,
   output        cfg_en2787,
   output        cfg_en2788,
   output        cfg_en2789,
   output        cfg_en2790,
   output        cfg_en2791,
   output        cfg_en2792,
   output        cfg_en2793,
   output        cfg_en2794,
   output        cfg_en2795,
   output        cfg_en2796,
   output        cfg_en2797,
   output        cfg_en2798,
   output        cfg_en2799,
   output        cfg_en2800,
   output        cfg_en2801,
   output        cfg_en2802,
   output        cfg_en2803,
   output        cfg_en2804,
   output        cfg_en2805,
   output        cfg_en2806,
   output        cfg_en2807,
   output        cfg_en2808,
   output        cfg_en2809,
   output        cfg_en2810,
   output        cfg_en2811,
   output        cfg_en2812,
   output        cfg_en2813,
   output        cfg_en2814,
   output        cfg_en2815,
   output        cfg_en2816,
   output        cfg_en2817,
   output        cfg_en2818,
   output        cfg_en2819,
   output        cfg_en2820,
   output        cfg_en2821,
   output        cfg_en2822,
   output        cfg_en2823,
   output        cfg_en2824,
   output        cfg_en2825,
   output        cfg_en2826,
   output        cfg_en2827,
   output        cfg_en2828,
   output        cfg_en2829,
   output        cfg_en2830,
   output        cfg_en2831,
   output        cfg_en2832,
   output        cfg_en2833,
   output        cfg_en2834,
   output        cfg_en2835,
   output        cfg_en2836,
   output        cfg_en2837,
   output        cfg_en2838,
   output        cfg_en2839,
   output        cfg_en2840,
   output        cfg_en2841,
   output        cfg_en2842,
   output        cfg_en2843,
   output        cfg_en2844,
   output        cfg_en2845,
   output        cfg_en2846,
   output        cfg_en2847,
   output        cfg_en2848,
   output        cfg_en2849,
   output        cfg_en2850,
   output        cfg_en2851,
   output        cfg_en2852,
   output        cfg_en2853,
   output        cfg_en2854,
   output        cfg_en2855,
   output        cfg_en2856,
   output        cfg_en2857,
   output        cfg_en2858,
   output        cfg_en2859,
   output        cfg_en2860,
   output        cfg_en2861,
   output        cfg_en2862,
   output        cfg_en2863,
   output        cfg_en2864,
   output        cfg_en2865,
   output        cfg_en2866,
   output        cfg_en2867,
   output        cfg_en2868,
   output        cfg_en2869,
   output        cfg_en2870,
   output        cfg_en2871,
   output        cfg_en2872,
   output        cfg_en2873,
   output        cfg_en2874,
   output        cfg_en2875,
   output        cfg_en2876,
   output        cfg_en2877,
   output        cfg_en2878,
   output        cfg_en2879,
   output        cfg_en2880,
   output        cfg_en2881,
   output        cfg_en2882,
   output        cfg_en2883,
   output        cfg_en2884,
   output        cfg_en2885,
   output        cfg_en2886,
   output        cfg_en2887,
   output        cfg_en2888,
   output        cfg_en2889,
   output        cfg_en2890,
   output        cfg_en2891,
   output        cfg_en2892,
   output        cfg_en2893,
   output        cfg_en2894,
   output        cfg_en2895,
   output        cfg_en2896,
   output        cfg_en2897,
   output        cfg_en2898,
   output        cfg_en2899,
   output        cfg_en2900,
   output        cfg_en2901,
   output        cfg_en2902,
   output        cfg_en2903,
   output        cfg_en2904,
   output        cfg_en2905,
   output        cfg_en2906,
   output        cfg_en2907,
   output        cfg_en2908,
   output        cfg_en2909,
   output        cfg_en2910,
   output        cfg_en2911,
   output        cfg_en2912,
   output        cfg_en2913,
   output        cfg_en2914,
   output        cfg_en2915,
   output        cfg_en2916,
   output        cfg_en2917,
   output        cfg_en2918,
   output        cfg_en2919,
   output        cfg_en2920,
   output        cfg_en2921,
   output        cfg_en2922,
   output        cfg_en2923,
   output        cfg_en2924,
   output        cfg_en2925,
   output        cfg_en2926,
   output        cfg_en2927,
   output        cfg_en2928,
   output        cfg_en2929,
   output        cfg_en2930,
   output        cfg_en2931,
   output        cfg_en2932,
   output        cfg_en2933,
   output        cfg_en2934,
   output        cfg_en2935,
   output        cfg_en2936,
   output        cfg_en2937,
   output        cfg_en2938,
   output        cfg_en2939,
   output        cfg_en2940,
   output        cfg_en2941,
   output        cfg_en2942,
   output        cfg_en2943,
   output        cfg_en2944,
   output        cfg_en2945,
   output        cfg_en2946,
   output        cfg_en2947,
   output        cfg_en2948,
   output        cfg_en2949,
   output        cfg_en2950,
   output        cfg_en2951,
   output        cfg_en2952,
   output        cfg_en2953,
   output        cfg_en2954,
   output        cfg_en2955,
   output        cfg_en2956,
   output        cfg_en2957,
   output        cfg_en2958,
   output        cfg_en2959,
   output        cfg_en2960,
   output        cfg_en2961,
   output        cfg_en2962,
   output        cfg_en2963,
   output        cfg_en2964,
   output        cfg_en2965,
   output        cfg_en2966,
   output        cfg_en2967,
   output        cfg_en2968,
   output        cfg_en2969,
   output        cfg_en2970,
   output        cfg_en2971,
   output        cfg_en2972,
   output        cfg_en2973,
   output        cfg_en2974,
   output        cfg_en2975,
   output        cfg_en2976,
   output        cfg_en2977,
   output        cfg_en2978,
   output        cfg_en2979,
   output        cfg_en2980,
   output        cfg_en2981,
   output        cfg_en2982,
   output        cfg_en2983,
   output        cfg_en2984,
   output        cfg_en2985,
   output        cfg_en2986,
   output        cfg_en2987,
   output        cfg_en2988,
   output        cfg_en2989,
   output        cfg_en2990,
   output        cfg_en2991,
   output        cfg_en2992,
   output        cfg_en2993,
   output        cfg_en2994,
   output        cfg_en2995,
   output        cfg_en2996,
   output        cfg_en2997,
   output        cfg_en2998,
   output        cfg_en2999,
   output        cfg_en3000,
   output        cfg_en3001,
   output        cfg_en3002,
   output        cfg_en3003,
   output        cfg_en3004,
   output        cfg_en3005,
   output        cfg_en3006,
   output        cfg_en3007,
   output        cfg_en3008,
   output        cfg_en3009,
   output        cfg_en3010,
   output        cfg_en3011,
   output        cfg_en3012,
   output        cfg_en3013,
   output        cfg_en3014,
   output        cfg_en3015,
   output        cfg_en3016,
   output        cfg_en3017,
   output        cfg_en3018,
   output        cfg_en3019,
   output        cfg_en3020,
   output        cfg_en3021,
   output        cfg_en3022,
   output        cfg_en3023,
   output        cfg_en3024,
   output        cfg_en3025,
   output        cfg_en3026,
   output        cfg_en3027,
   output        cfg_en3028,
   output        cfg_en3029,
   output        cfg_en3030,
   output        cfg_en3031,
   output        cfg_en3032,
   output        cfg_en3033,
   output        cfg_en3034,
   output        cfg_en3035,
   output        cfg_en3036,
   output        cfg_en3037,
   output        cfg_en3038,
   output        cfg_en3039,
   output        cfg_en3040,
   output        cfg_en3041,
   output        cfg_en3042,
   output        cfg_en3043,
   output        cfg_en3044,
   output        cfg_en3045,
   output        cfg_en3046,
   output        cfg_en3047,
   output        cfg_en3048,
   output        cfg_en3049,
   output        cfg_en3050,
   output        cfg_en3051,
   output        cfg_en3052,
   output        cfg_en3053,
   output        cfg_en3054,
   output        cfg_en3055,
   output        cfg_en3056,
   output        cfg_en3057,
   output        cfg_en3058,
   output        cfg_en3059,
   output        cfg_en3060,
   output        cfg_en3061,
   output        cfg_en3062,
   output        cfg_en3063,
   output        cfg_en3064,
   output        cfg_en3065,
   output        cfg_en3066,
   output        cfg_en3067,
   output        cfg_en3068,
   output        cfg_en3069,
   output        cfg_en3070,
   output        cfg_en3071,
   output        cfg_en3072,
   output        cfg_en3073,
   output        cfg_en3074,
   output        cfg_en3075,
   output        cfg_en3076,
   output        cfg_en3077,
   output        cfg_en3078,
   output        cfg_en3079,
   output        cfg_en3080,
   output        cfg_en3081,
   output        cfg_en3082,
   output        cfg_en3083,
   output        cfg_en3084,
   output        cfg_en3085,
   output        cfg_en3086,
   output        cfg_en3087,
   output        cfg_en3088,
   output        cfg_en3089,
   output        cfg_en3090,
   output        cfg_en3091,
   output        cfg_en3092,
   output        cfg_en3093,
   output        cfg_en3094,
   output        cfg_en3095,
   output        cfg_en3096,
   output        cfg_en3097,
   output        cfg_en3098,
   output        cfg_en3099,
   output        cfg_en3100,
   output        cfg_en3101,
   output        cfg_en3102,
   output        cfg_en3103,
   output        cfg_en3104,
   output        cfg_en3105,
   output        cfg_en3106,
   output        cfg_en3107,
   output        cfg_en3108,
   output        cfg_en3109,
   output        cfg_en3110,
   output        cfg_en3111,
   output        cfg_en3112,
   output        cfg_en3113,
   output        cfg_en3114,
   output        cfg_en3115,
   output        cfg_en3116,
   output        cfg_en3117,
   output        cfg_en3118,
   output        cfg_en3119,
   output        cfg_en3120,
   output        cfg_en3121,
   output        cfg_en3122,
   output        cfg_en3123,
   output        cfg_en3124,
   output        cfg_en3125,
   output        cfg_en3126,
   output        cfg_en3127,
   output        cfg_en3128,
   output        cfg_en3129,
   output        cfg_en3130,
   output        cfg_en3131,
   output        cfg_en3132,
   output        cfg_en3133,
   output        cfg_en3134,
   output        cfg_en3135,
   output        cfg_en3136,
   output        cfg_en3137,
   output        cfg_en3138,
   output        cfg_en3139,
   output        cfg_en3140,
   output        cfg_en3141,
   output        cfg_en3142,
   output        cfg_en3143,
   output        cfg_en3144,
   output        cfg_en3145,
   output        cfg_en3146,
   output        cfg_en3147,
   output        cfg_en3148,
   output        cfg_en3149,
   output        cfg_en3150,
   output        cfg_en3151,
   output        cfg_en3152,
   output        cfg_en3153,
   output        cfg_en3154,
   output        cfg_en3155,
   output        cfg_en3156,
   output        cfg_en3157,
   output        cfg_en3158,
   output        cfg_en3159,
   output        cfg_en3160,
   output        cfg_en3161,
   output        cfg_en3162,
   output        cfg_en3163,
   output        cfg_en3164,
   output        cfg_en3165,
   output        cfg_en3166,
   output        cfg_en3167,
   output        cfg_en3168,
   output        cfg_en3169,
   output        cfg_en3170,
   output        cfg_en3171,
   output        cfg_en3172,
   output        cfg_en3173,
   output        cfg_en3174,
   output        cfg_en3175,
   output        cfg_en3176,
   output        cfg_en3177,
   output        cfg_en3178,
   output        cfg_en3179,
   output        cfg_en3180,
   output        cfg_en3181,
   output        cfg_en3182,
   output        cfg_en3183,
   output        cfg_en3184,
   output        cfg_en3185,
   output        cfg_en3186,
   output        cfg_en3187,
   output        cfg_en3188,
   output        cfg_en3189,
   output        cfg_en3190,
   output        cfg_en3191,
   output        cfg_en3192,
   output        cfg_en3193,
   output        cfg_en3194,
   output        cfg_en3195,
   output        cfg_en3196,
   output        cfg_en3197,
   output        cfg_en3198,
   output        cfg_en3199,
   output        cfg_en3200,
   output        cfg_en3201,
   output        cfg_en3202,
   output        cfg_en3203,
   output        cfg_en3204,
   output        cfg_en3205,
   output        cfg_en3206,
   output        cfg_en3207,
   output        cfg_en3208,
   output        cfg_en3209,
   output        cfg_en3210,
   output        cfg_en3211,
   output        cfg_en3212,
   output        cfg_en3213,
   output        cfg_en3214,
   output        cfg_en3215,
   output        cfg_en3216,
   output        cfg_en3217,
   output        cfg_en3218,
   output        cfg_en3219,
   output        cfg_en3220,
   output        cfg_en3221,
   output        cfg_en3222,
   output        cfg_en3223,
   output        cfg_en3224,
   output        cfg_en3225,
   output        cfg_en3226,
   output        cfg_en3227,
   output        cfg_en3228,
   output        cfg_en3229,
   output        cfg_en3230,
   output        cfg_en3231,
   output        cfg_en3232,
   output        cfg_en3233,
   output        cfg_en3234,
   output        cfg_en3235,
   output        cfg_en3236,
   output        cfg_en3237,
   output        cfg_en3238,
   output        cfg_en3239,
   output        cfg_en3240,
   output        cfg_en3241,
   output        cfg_en3242,
   output        cfg_en3243,
   output        cfg_en3244,
   output        cfg_en3245,
   output        cfg_en3246,
   output        cfg_en3247,
   output        cfg_en3248,
   output        cfg_en3249,
   output        cfg_en3250,
   output        cfg_en3251,
   output        cfg_en3252,
   output        cfg_en3253,
   output        cfg_en3254,
   output        cfg_en3255,
   output        cfg_en3256,
   output        cfg_en3257,
   output        cfg_en3258,
   output        cfg_en3259,
   output        cfg_en3260,
   output        cfg_en3261,
   output        cfg_en3262,
   output        cfg_en3263,
   output        cfg_en3264,
   output        cfg_en3265,
   output        cfg_en3266,
   output        cfg_en3267,
   output        cfg_en3268,
   output        cfg_en3269,
   output        cfg_en3270,
   output        cfg_en3271,
   output        cfg_en3272,
   output        cfg_en3273,
   output        cfg_en3274,
   output        cfg_en3275,
   output        cfg_en3276,
   output        cfg_en3277,
   output        cfg_en3278,
   output        cfg_en3279,
   output        cfg_en3280,
   output        cfg_en3281,
   output        cfg_en3282,
   output        cfg_en3283,
   output        cfg_en3284,
   output        cfg_en3285,
   output        cfg_en3286,
   output        cfg_en3287,
   output        cfg_en3288,
   output        cfg_en3289,
   output        cfg_en3290,
   output        cfg_en3291,
   output        cfg_en3292,
   output        cfg_en3293,
   output        cfg_en3294,
   output        cfg_en3295,
   output        cfg_en3296,
   output        cfg_en3297,
   output        cfg_en3298,
   output        cfg_en3299,
   output        cfg_en3300,
   output        cfg_en3301,
   output        cfg_en3302,
   output        cfg_en3303,
   output        cfg_en3304,
   output        cfg_en3305,
   output        cfg_en3306,
   output        cfg_en3307,
   output        cfg_en3308,
   output        cfg_en3309,
   output        cfg_en3310,
   output        cfg_en3311,
   output        cfg_en3312,
   output        cfg_en3313,
   output        cfg_en3314,
   output        cfg_en3315,
   output        cfg_en3316,
   output        cfg_en3317,
   output        cfg_en3318,
   output        cfg_en3319,
   output        cfg_en3320,
   output        cfg_en3321,
   output        cfg_en3322,
   output        cfg_en3323,
   output        cfg_en3324,
   output        cfg_en3325,
   output        cfg_en3326,
   output        cfg_en3327,
   output        cfg_en3328,
   output        cfg_en3329,
   output        cfg_en3330,
   output        cfg_en3331,
   output        cfg_en3332,
   output        cfg_en3333,
   output        cfg_en3334,
   output        cfg_en3335,
   output        cfg_en3336,
   output        cfg_en3337,
   output        cfg_en3338,
   output        cfg_en3339,
   output        cfg_en3340,
   output        cfg_en3341,
   output        cfg_en3342,
   output        cfg_en3343,
   output        cfg_en3344,
   output        cfg_en3345,
   output        cfg_en3346,
   output        cfg_en3347,
   output        cfg_en3348,
   output        cfg_en3349,
   output        cfg_en3350,
   output        cfg_en3351,
   output        cfg_en3352,
   output        cfg_en3353,
   output        cfg_en3354,
   output        cfg_en3355,
   output        cfg_en3356,
   output        cfg_en3357,
   output        cfg_en3358,
   output        cfg_en3359,
   output        cfg_en3360,
   output        cfg_en3361,
   output        cfg_en3362,
   output        cfg_en3363,
   output        cfg_en3364,
   output        cfg_en3365,
   output        cfg_en3366,
   output        cfg_en3367,
   output        cfg_en3368,
   output        cfg_en3369,
   output        cfg_en3370,
   output        cfg_en3371,
   output        cfg_en3372,
   output        cfg_en3373,
   output        cfg_en3374,
   output        cfg_en3375,
   output        cfg_en3376,
   output        cfg_en3377,
   output        cfg_en3378,
   output        cfg_en3379,
   output        cfg_en3380,
   output        cfg_en3381,
   output        cfg_en3382,
   output        cfg_en3383,
   output        cfg_en3384,
   output        cfg_en3385,
   output        cfg_en3386,
   output        cfg_en3387,
   output        cfg_en3388,
   output        cfg_en3389,
   output        cfg_en3390,
   output        cfg_en3391,
   output        cfg_en3392,
   output        cfg_en3393,
   output        cfg_en3394,
   output        cfg_en3395,
   output        cfg_en3396,
   output        cfg_en3397,
   output        cfg_en3398,
   output        cfg_en3399,
   output        cfg_en3400,
   output        cfg_en3401,
   output        cfg_en3402,
   output        cfg_en3403,
   output        cfg_en3404,
   output        cfg_en3405,
   output        cfg_en3406,
   output        cfg_en3407,
   output        cfg_en3408,
   output        cfg_en3409,
   output        cfg_en3410,
   output        cfg_en3411,
   output        cfg_en3412,
   output        cfg_en3413,
   output        cfg_en3414,
   output        cfg_en3415,
   output        cfg_en3416,
   output        cfg_en3417,
   output        cfg_en3418,
   output        cfg_en3419,
   output        cfg_en3420,
   output        cfg_en3421,
   output        cfg_en3422,
   output        cfg_en3423,
   output        cfg_en3424,
   output        cfg_en3425,
   output        cfg_en3426,
   output        cfg_en3427,
   output        cfg_en3428,
   output        cfg_en3429,
   output        cfg_en3430,
   output        cfg_en3431,
   output        cfg_en3432,
   output        cfg_en3433,
   output        cfg_en3434,
   output        cfg_en3435,
   output        cfg_en3436,
   output        cfg_en3437,
   output        cfg_en3438,
   output        cfg_en3439,
   output        cfg_en3440,
   output        cfg_en3441,
   output        cfg_en3442,
   output        cfg_en3443,
   output        cfg_en3444,
   output        cfg_en3445,
   output        cfg_en3446,
   output        cfg_en3447,
   output        cfg_en3448,
   output        cfg_en3449,
   output        cfg_en3450,
   output        cfg_en3451,
   output        cfg_en3452,
   output        cfg_en3453,
   output        cfg_en3454,
   output        cfg_en3455,
   output        cfg_en3456,
   output        cfg_en3457,
   output        cfg_en3458,
   output        cfg_en3459,
   output        cfg_en3460,
   output        cfg_en3461,
   output        cfg_en3462,
   output        cfg_en3463,
   output        cfg_en3464,
   output        cfg_en3465,
   output        cfg_en3466,
   output        cfg_en3467,
   output        cfg_en3468,
   output        cfg_en3469,
   output        cfg_en3470,
   output        cfg_en3471,
   output        cfg_en3472,
   output        cfg_en3473,
   output        cfg_en3474,
   output        cfg_en3475,
   output        cfg_en3476,
   output        cfg_en3477,
   output        cfg_en3478,
   output        cfg_en3479,
   output        cfg_en3480,
   output        cfg_en3481,
   output        cfg_en3482,
   output        cfg_en3483,
   output        cfg_en3484,
   output        cfg_en3485,
   output        cfg_en3486,
   output        cfg_en3487,
   output        cfg_en3488,
   output        cfg_en3489,
   output        cfg_en3490,
   output        cfg_en3491,
   output        cfg_en3492,
   output        cfg_en3493,
   output        cfg_en3494,
   output        cfg_en3495,
   output        cfg_en3496,
   output        cfg_en3497,
   output        cfg_en3498,
   output        cfg_en3499,
   output        cfg_en3500,
   output        cfg_en3501,
   output        cfg_en3502,
   output        cfg_en3503,
   output        cfg_en3504,
   output        cfg_en3505,
   output        cfg_en3506,
   output        cfg_en3507,
   output        cfg_en3508,
   output        cfg_en3509,
   output        cfg_en3510,
   output        cfg_en3511,
   output        cfg_en3512,
   output        cfg_en3513,
   output        cfg_en3514,
   output        cfg_en3515,
   output        cfg_en3516,
   output        cfg_en3517,
   output        cfg_en3518,
   output        cfg_en3519,
   output        cfg_en3520,
   output        cfg_en3521,
   output        cfg_en3522,
   output        cfg_en3523,
   output        cfg_en3524,
   output        cfg_en3525,
   output        cfg_en3526,
   output        cfg_en3527,
   output        cfg_en3528,
   output        cfg_en3529,
   output        cfg_en3530,
   output        cfg_en3531,
   output        cfg_en3532,
   output        cfg_en3533,
   output        cfg_en3534,
   output        cfg_en3535,
   output        cfg_en3536,
   output        cfg_en3537,
   output        cfg_en3538,
   output        cfg_en3539,
   output        cfg_en3540,
   output        cfg_en3541,
   output        cfg_en3542,
   output        cfg_en3543,
   output        cfg_en3544,
   output        cfg_en3545,
   output        cfg_en3546,
   output        cfg_en3547,
   output        cfg_en3548,
   output        cfg_en3549,
   output        cfg_en3550,
   output        cfg_en3551,
   output        cfg_en3552,
   output        cfg_en3553,
   output        cfg_en3554,
   output        cfg_en3555,
   output        cfg_en3556,
   output        cfg_en3557,
   output        cfg_en3558,
   output        cfg_en3559,
   output        cfg_en3560,
   output        cfg_en3561,
   output        cfg_en3562,
   output        cfg_en3563,
   output        cfg_en3564,
   output        cfg_en3565,
   output        cfg_en3566,
   output        cfg_en3567,
   output        cfg_en3568,
   output        cfg_en3569,
   output        cfg_en3570,
   output        cfg_en3571,
   output        cfg_en3572,
   output        cfg_en3573,
   output        cfg_en3574,
   output        cfg_en3575,
   output        cfg_en3576,
   output        cfg_en3577,
   output        cfg_en3578,
   output        cfg_en3579,
   output        cfg_en3580,
   output        cfg_en3581,
   output        cfg_en3582,
   output        cfg_en3583,
   output        cfg_en3584,
   output        cfg_en3585,
   output        cfg_en3586,
   output        cfg_en3587,
   output        cfg_en3588,
   output        cfg_en3589,
   output        cfg_en3590,
   output        cfg_en3591,
   output        cfg_en3592,
   output        cfg_en3593,
   output        cfg_en3594,
   output        cfg_en3595,
   output        cfg_en3596,
   output        cfg_en3597,
   output        cfg_en3598,
   output        cfg_en3599,
   output        cfg_en3600,
   output        cfg_en3601,
   output        cfg_en3602,
   output        cfg_en3603,
   output        cfg_en3604,
   output        cfg_en3605,
   output        cfg_en3606,
   output        cfg_en3607,
   output        cfg_en3608,
   output        cfg_en3609,
   output        cfg_en3610,
   output        cfg_en3611,
   output        cfg_en3612,
   output        cfg_en3613,
   output        cfg_en3614,
   output        cfg_en3615,
   output        cfg_en3616,
   output        cfg_en3617,
   output        cfg_en3618,
   output        cfg_en3619,
   output        cfg_en3620,
   output        cfg_en3621,
   output        cfg_en3622,
   output        cfg_en3623,
   output        cfg_en3624,
   output        cfg_en3625,
   output        cfg_en3626,
   output        cfg_en3627,
   output        cfg_en3628,
   output        cfg_en3629,
   output        cfg_en3630,
   output        cfg_en3631,
   output        cfg_en3632,
   output        cfg_en3633,
   output        cfg_en3634,
   output        cfg_en3635,
   output        cfg_en3636,
   output        cfg_en3637,
   output        cfg_en3638,
   output        cfg_en3639,
   output        cfg_en3640,
   output        cfg_en3641,
   output        cfg_en3642,
   output        cfg_en3643,
   output        cfg_en3644,
   output        cfg_en3645,
   output        cfg_en3646,
   output        cfg_en3647,
   output        cfg_en3648,
   output        cfg_en3649,
   output        cfg_en3650,
   output        cfg_en3651,
   output        cfg_en3652,
   output        cfg_en3653,
   output        cfg_en3654,
   output        cfg_en3655,
   output        cfg_en3656,
   output        cfg_en3657,
   output        cfg_en3658,
   output        cfg_en3659,
   output        cfg_en3660,
   output        cfg_en3661,
   output        cfg_en3662,
   output        cfg_en3663,
   output        cfg_en3664,
   output        cfg_en3665,
   output        cfg_en3666,
   output        cfg_en3667,
   output        cfg_en3668,
   output        cfg_en3669,
   output        cfg_en3670,
   output        cfg_en3671,
   output        cfg_en3672,
   output        cfg_en3673,
   output        cfg_en3674,
   output        cfg_en3675,
   output        cfg_en3676,
   output        cfg_en3677,
   output        cfg_en3678,
   output        cfg_en3679,
   output        cfg_en3680,
   output        cfg_en3681,
   output        cfg_en3682,
   output        cfg_en3683,
   output        cfg_en3684,
   output        cfg_en3685,
   output        cfg_en3686,
   output        cfg_en3687,
   output        cfg_en3688,
   output        cfg_en3689,
   output        cfg_en3690,
   output        cfg_en3691,
   output        cfg_en3692,
   output        cfg_en3693,
   output        cfg_en3694,
   output        cfg_en3695,
   output        cfg_en3696,
   output        cfg_en3697,
   output        cfg_en3698,
   output        cfg_en3699,
   output        cfg_en3700,
   output        cfg_en3701,
   output        cfg_en3702,
   output        cfg_en3703,
   output        cfg_en3704,
   output        cfg_en3705,
   output        cfg_en3706,
   output        cfg_en3707,
   output        cfg_en3708,
   output        cfg_en3709,
   output        cfg_en3710,
   output        cfg_en3711,
   output        cfg_en3712,
   output        cfg_en3713,
   output        cfg_en3714,
   output        cfg_en3715,
   output        cfg_en3716,
   output        cfg_en3717,
   output        cfg_en3718,
   output        cfg_en3719,
   output        cfg_en3720,
   output        cfg_en3721,
   output        cfg_en3722,
   output        cfg_en3723,
   output        cfg_en3724,
   output        cfg_en3725,
   output        cfg_en3726,
   output        cfg_en3727,
   output        cfg_en3728,
   output        cfg_en3729,
   output        cfg_en3730,
   output        cfg_en3731,
   output        cfg_en3732,
   output        cfg_en3733,
   output        cfg_en3734,
   output        cfg_en3735,
   output        cfg_en3736,
   output        cfg_en3737,
   output        cfg_en3738,
   output        cfg_en3739,
   output        cfg_en3740,
   output        cfg_en3741,
   output        cfg_en3742,
   output        cfg_en3743,
   output        cfg_en3744,
   output        cfg_en3745,
   output        cfg_en3746,
   output        cfg_en3747,
   output        cfg_en3748,
   output        cfg_en3749,
   output        cfg_en3750,
   output        cfg_en3751,
   output        cfg_en3752,
   output        cfg_en3753,
   output        cfg_en3754,
   output        cfg_en3755,
   output        cfg_en3756,
   output        cfg_en3757,
   output        cfg_en3758,
   output        cfg_en3759,
   output        cfg_en3760,
   output        cfg_en3761,
   output        cfg_en3762,
   output        cfg_en3763,
   output        cfg_en3764,
   output        cfg_en3765,
   output        cfg_en3766,
   output        cfg_en3767,
   output        cfg_en3768,
   output        cfg_en3769,
   output        cfg_en3770,
   output        cfg_en3771,
   output        cfg_en3772,
   output        cfg_en3773,
   output        cfg_en3774,
   output        cfg_en3775,
   output        cfg_en3776,
   output        cfg_en3777,
   output        cfg_en3778,
   output        cfg_en3779,
   output        cfg_en3780,
   output        cfg_en3781,
   output        cfg_en3782,
   output        cfg_en3783,
   output        cfg_en3784,
   output        cfg_en3785,
   output        cfg_en3786,
   output        cfg_en3787,
   output        cfg_en3788,
   output        cfg_en3789,
   output        cfg_en3790,
   output        cfg_en3791,
   output        cfg_en3792,
   output        cfg_en3793,
   output        cfg_en3794,
   output        cfg_en3795,
   output        cfg_en3796,
   output        cfg_en3797,
   output        cfg_en3798,
   output        cfg_en3799,
   output        cfg_en3800,
   output        cfg_en3801,
   output        cfg_en3802,
   output        cfg_en3803,
   output        cfg_en3804,
   output        cfg_en3805,
   output        cfg_en3806,
   output        cfg_en3807,
   output        cfg_en3808,
   output        cfg_en3809,
   output        cfg_en3810,
   output        cfg_en3811,
   output        cfg_en3812,
   output        cfg_en3813,
   output        cfg_en3814,
   output        cfg_en3815,
   output        cfg_en3816,
   output        cfg_en3817,
   output        cfg_en3818,
   output        cfg_en3819,
   output        cfg_en3820,
   output        cfg_en3821,
   output        cfg_en3822,
   output        cfg_en3823,
   output        cfg_en3824,
   output        cfg_en3825,
   output        cfg_en3826,
   output        cfg_en3827,
   output        cfg_en3828,
   output        cfg_en3829,
   output        cfg_en3830,
   output        cfg_en3831,
   output        cfg_en3832,
   output        cfg_en3833,
   output        cfg_en3834,
   output        cfg_en3835,
   output        cfg_en3836,
   output        cfg_en3837,
   output        cfg_en3838,
   output        cfg_en3839,
   output        cfg_en3840,
   output        cfg_en3841,
   output        cfg_en3842,
   output        cfg_en3843,
   output        cfg_en3844,
   output        cfg_en3845,
   output        cfg_en3846,
   output        cfg_en3847,
   output        cfg_en3848,
   output        cfg_en3849,
   output        cfg_en3850,
   output        cfg_en3851,
   output        cfg_en3852,
   output        cfg_en3853,
   output        cfg_en3854,
   output        cfg_en3855,
   output        cfg_en3856,
   output        cfg_en3857,
   output        cfg_en3858,
   output        cfg_en3859,
   output        cfg_en3860,
   output        cfg_en3861,
   output        cfg_en3862,
   output        cfg_en3863,
   output        cfg_en3864,
   output        cfg_en3865,
   output        cfg_en3866,
   output        cfg_en3867,
   output        cfg_en3868,
   output        cfg_en3869,
   output        cfg_en3870,
   output        cfg_en3871,
   output        cfg_en3872,
   output        cfg_en3873,
   output        cfg_en3874,
   output        cfg_en3875,
   output        cfg_en3876,
   output        cfg_en3877,
   output        cfg_en3878,
   output        cfg_en3879,
   output        cfg_en3880,
   output        cfg_en3881,
   output        cfg_en3882,
   output        cfg_en3883,
   output        cfg_en3884,
   output        cfg_en3885,
   output        cfg_en3886,
   output        cfg_en3887,
   output        cfg_en3888,
   output        cfg_en3889,
   output        cfg_en3890,
   output        cfg_en3891,
   output        cfg_en3892,
   output        cfg_en3893,
   output        cfg_en3894,
   output        cfg_en3895,
   output        cfg_en3896,
   output        cfg_en3897,
   output        cfg_en3898,
   output        cfg_en3899,
   output        cfg_en3900,
   output        cfg_en3901,
   output        cfg_en3902,
   output        cfg_en3903,
   output        cfg_en3904,
   output        cfg_en3905,
   output        cfg_en3906,
   output        cfg_en3907,
   output        cfg_en3908,
   output        cfg_en3909,
   output        cfg_en3910,
   output        cfg_en3911,
   output        cfg_en3912,
   output        cfg_en3913,
   output        cfg_en3914,
   output        cfg_en3915,
   output        cfg_en3916,
   output        cfg_en3917,
   output        cfg_en3918,
   output        cfg_en3919,
   output        cfg_en3920,
   output        cfg_en3921,
   output        cfg_en3922,
   output        cfg_en3923,
   output        cfg_en3924,
   output        cfg_en3925,
   output        cfg_en3926,
   output        cfg_en3927,
   output        cfg_en3928,
   output        cfg_en3929,
   output        cfg_en3930,
   output        cfg_en3931,
   output        cfg_en3932,
   output        cfg_en3933,
   output        cfg_en3934,
   output        cfg_en3935,
   output        cfg_en3936,
   output        cfg_en3937,
   output        cfg_en3938,
   output        cfg_en3939,
   output        cfg_en3940,
   output        cfg_en3941,
   output        cfg_en3942,
   output        cfg_en3943,
   output        cfg_en3944,
   output        cfg_en3945,
   output        cfg_en3946,
   output        cfg_en3947,
   output        cfg_en3948,
   output        cfg_en3949,
   output        cfg_en3950,
   output        cfg_en3951,
   output        cfg_en3952,
   output        cfg_en3953,
   output        cfg_en3954,
   output        cfg_en3955,
   output        cfg_en3956,
   output        cfg_en3957,
   output        cfg_en3958,
   output        cfg_en3959,
   output        cfg_en3960,
   output        cfg_en3961,
   output        cfg_en3962,
   output        cfg_en3963,
   output        cfg_en3964,
   output        cfg_en3965,
   output        cfg_en3966,
   output        cfg_en3967,
   output        cfg_en3968,
   output        cfg_en3969,
   output        cfg_en3970,
   output        cfg_en3971,
   output        cfg_en3972,
   output        cfg_en3973,
   output        cfg_en3974,
   output        cfg_en3975,
   output        cfg_en3976,
   output        cfg_en3977,
   output        cfg_en3978,
   output        cfg_en3979,
   output        cfg_en3980,
   output        cfg_en3981,
   output        cfg_en3982,
   output        cfg_en3983,
   output        cfg_en3984,
   output        cfg_en3985,
   output        cfg_en3986,
   output        cfg_en3987,
   output        cfg_en3988,
   output        cfg_en3989,
   output        cfg_en3990,
   output        cfg_en3991,
   output        cfg_en3992,
   output        cfg_en3993,
   output        cfg_en3994,
   output        cfg_en3995,
   output        cfg_en3996,
   output        cfg_en3997,
   output        cfg_en3998,
   output        cfg_en3999,
   output        cfg_en4000,
   output        cfg_en4001,
   output        cfg_en4002,
   output        cfg_en4003,
   output        cfg_en4004,
   output        cfg_en4005,
   output        cfg_en4006,
   output        cfg_en4007,
   output        cfg_en4008,
   output        cfg_en4009,
   output        cfg_en4010,
   output        cfg_en4011,
   output        cfg_en4012,
   output        cfg_en4013,
   output        cfg_en4014,
   output        cfg_en4015,
   output        cfg_en4016,
   output        cfg_en4017,
   output        cfg_en4018,
   output        cfg_en4019,
   output        cfg_en4020,
   output        cfg_en4021,
   output        cfg_en4022,
   output        cfg_en4023,
   output        cfg_en4024,
   output        cfg_en4025,
   output        cfg_en4026,
   output        cfg_en4027,
   output        cfg_en4028,
   output        cfg_en4029,
   output        cfg_en4030,
   output        cfg_en4031,
   output        cfg_en4032,
   output        cfg_en4033,
   output        cfg_en4034,
   output        cfg_en4035,
   output        cfg_en4036,
   output        cfg_en4037,
   output        cfg_en4038,
   output        cfg_en4039,
   output        cfg_en4040,
   output        cfg_en4041,
   output        cfg_en4042,
   output        cfg_en4043,
   output        cfg_en4044,
   output        cfg_en4045,
   output        cfg_en4046,
   output        cfg_en4047,
   output        cfg_en4048,
   output        cfg_en4049,
   output        cfg_en4050,
   output        cfg_en4051,
   output        cfg_en4052,
   output        cfg_en4053,
   output        cfg_en4054,
   output        cfg_en4055,
   output        cfg_en4056,
   output        cfg_en4057,
   output        cfg_en4058,
   output        cfg_en4059,
   output        cfg_en4060,
   output        cfg_en4061,
   output        cfg_en4062,
   output        cfg_en4063,
   output        cfg_en4064,
   output        cfg_en4065,
   output        cfg_en4066,
   output        cfg_en4067,
   output        cfg_en4068,
   output        cfg_en4069,
   output        cfg_en4070,
   output        cfg_en4071,
   output        cfg_en4072,
   output        cfg_en4073,
   output        cfg_en4074,
   output        cfg_en4075,
   output        cfg_en4076,
   output        cfg_en4077,
   output        cfg_en4078,
   output        cfg_en4079,
   output        cfg_en4080,
   output        cfg_en4081,
   output        cfg_en4082,
   output        cfg_en4083,
   output        cfg_en4084,
   output        cfg_en4085,
   output        cfg_en4086,
   output        cfg_en4087,
   output        cfg_en4088,
   output        cfg_en4089,
   output        cfg_en4090,
   output        cfg_en4091,
   output        cfg_en4092,
   output        cfg_en4093,
   output        cfg_en4094,
   output        cfg_en4095,
   output        tc_cfg_en,
   output        cc_cfg_en0,
   output        cc_cfg_en1,
   output        cc_cfg_en2,
   output        cc_cfg_en3,
   output        cfg_din0,
   output        cfg_din1,
   output        cfg_din2,
   output        cfg_din3,
   output        cfg_din4,
   output        cfg_din5,
   output        cfg_din6,
   output        cfg_din7,
   output        cfg_din8,
   output        cfg_din9,
   output        cfg_din10,
   output        cfg_din11,
   output        cfg_din12,
   output        cfg_din13,
   output        cfg_din14,
   output        cfg_din15,
   output        cfg_din16,
   output        cfg_din17,
   output        cfg_din18,
   output        cfg_din19,
   output        cfg_din20,
   output        cfg_din21,
   output        cfg_din22,
   output        cfg_din23,
   output        cfg_din24,
   output        cfg_din25,
   output        cfg_din26,
   output        cfg_din27,
   output        cfg_din28,
   output        cfg_din29,
   output        cfg_din30,
   output        cfg_din31,
   output        cfg_din32,
   output        cfg_din33,
   output        cfg_din34,
   output        cfg_din35,
   output        cfg_din36,
   output        cfg_din37,
   output        cfg_din38,
   output        cfg_din39,
   output        cfg_din40,
   output        cfg_din41,
   output        cfg_din42,
   output        cfg_din43,
   output        cfg_din44,
   output        cfg_din45,
   output        cfg_din46,
   output        cfg_din47,
   output        cfg_din48,
   output        cfg_din49,
   output        cfg_din50,
   output        cfg_din51,
   output        cfg_din52,
   output        cfg_din53,
   output        cfg_din54,
   output        cfg_din55,
   output        cfg_din56,
   output        cfg_din57,
   output        cfg_din58,
   output        cfg_din59,
   output        cfg_din60,
   output        cfg_din61,
   output        cfg_din62,
   output        cfg_din63,
   output        cfg_din64,
   output        cfg_din65,
   output        cfg_din66,
   output        cfg_din67,
   output        cfg_din68,
   output        cfg_din69,
   output        cfg_din70,
   output        cfg_din71,
   output        cfg_din72,
   output        cfg_din73,
   output        cfg_din74,
   output        cfg_din75,
   output        cfg_din76,
   output        cfg_din77,
   output        cfg_din78,
   output        cfg_din79,
   output        cfg_din80,
   output        cfg_din81,
   output        cfg_din82,
   output        cfg_din83,
   output        cfg_din84,
   output        cfg_din85,
   output        cfg_din86,
   output        cfg_din87,
   output        cfg_din88,
   output        cfg_din89,
   output        cfg_din90,
   output        cfg_din91,
   output        cfg_din92,
   output        cfg_din93,
   output        cfg_din94,
   output        cfg_din95,
   output        cfg_din96,
   output        cfg_din97,
   output        cfg_din98,
   output        cfg_din99,
   output        cfg_din100,
   output        cfg_din101,
   output        cfg_din102,
   output        cfg_din103,
   output        cfg_din104,
   output        cfg_din105,
   output        cfg_din106,
   output        cfg_din107,
   output        cfg_din108,
   output        cfg_din109,
   output        cfg_din110,
   output        cfg_din111,
   output        cfg_din112,
   output        cfg_din113,
   output        cfg_din114,
   output        cfg_din115,
   output        cfg_din116,
   output        cfg_din117,
   output        cfg_din118,
   output        cfg_din119,
   output        cfg_din120,
   output        cfg_din121,
   output        cfg_din122,
   output        cfg_din123,
   output        cfg_din124,
   output        cfg_din125,
   output        cfg_din126,
   output        cfg_din127,
   output        cfg_din128,
   output        cfg_din129,
   output        cfg_din130,
   output        cfg_din131,
   output        cfg_din132,
   output        cfg_din133,
   output        cfg_din134,
   output        cfg_din135,
   output        cfg_din136,
   output        cfg_din137,
   output        cfg_din138,
   output        cfg_din139,
   output        cfg_din140,
   output        cfg_din141,
   output        cfg_din142,
   output        cfg_din143,
   output        cfg_din144,
   output        cfg_din145,
   output        cfg_din146,
   output        cfg_din147,
   output        cfg_din148,
   output        cfg_din149,
   output        cfg_din150,
   output        cfg_din151,
   output        cfg_din152,
   output        cfg_din153,
   output        cfg_din154,
   output        cfg_din155,
   output        cfg_din156,
   output        cfg_din157,
   output        cfg_din158,
   output        cfg_din159,
   output        cfg_din160,
   output        cfg_din161,
   output        cfg_din162,
   output        cfg_din163,
   output        cfg_din164,
   output        cfg_din165,
   output        cfg_din166,
   output        cfg_din167,
   output        cfg_din168,
   output        cfg_din169,
   output        cfg_din170,
   output        cfg_din171,
   output        cfg_din172,
   output        cfg_din173,
   output        cfg_din174,
   output        cfg_din175,
   output        cfg_din176,
   output        cfg_din177,
   output        cfg_din178,
   output        cfg_din179,
   output        cfg_din180,
   output        cfg_din181,
   output        cfg_din182,
   output        cfg_din183,
   output        cfg_din184,
   output        cfg_din185,
   output        cfg_din186,
   output        cfg_din187,
   output        cfg_din188,
   output        cfg_din189,
   output        cfg_din190,
   output        cfg_din191,
   output        cfg_din192,
   output        cfg_din193,
   output        cfg_din194,
   output        cfg_din195,
   output        cfg_din196,
   output        cfg_din197,
   output        cfg_din198,
   output        cfg_din199,
   output        cfg_din200,
   output        cfg_din201,
   output        cfg_din202,
   output        cfg_din203,
   output        cfg_din204,
   output        cfg_din205,
   output        cfg_din206,
   output        cfg_din207,
   output        cfg_din208,
   output        cfg_din209,
   output        cfg_din210,
   output        cfg_din211,
   output        cfg_din212,
   output        cfg_din213,
   output        cfg_din214,
   output        cfg_din215,
   output        cfg_din216,
   output        cfg_din217,
   output        cfg_din218,
   output        cfg_din219,
   output        cfg_din220,
   output        cfg_din221,
   output        cfg_din222,
   output        cfg_din223,
   output        cfg_din224,
   output        cfg_din225,
   output        cfg_din226,
   output        cfg_din227,
   output        cfg_din228,
   output        cfg_din229,
   output        cfg_din230,
   output        cfg_din231,
   output        cfg_din232,
   output        cfg_din233,
   output        cfg_din234,
   output        cfg_din235,
   output        cfg_din236,
   output        cfg_din237,
   output        cfg_din238,
   output        cfg_din239,
   output        cfg_din240,
   output        cfg_din241,
   output        cfg_din242,
   output        cfg_din243,
   output        cfg_din244,
   output        cfg_din245,
   output        cfg_din246,
   output        cfg_din247,
   output        cfg_din248,
   output        cfg_din249,
   output        cfg_din250,
   output        cfg_din251,
   output        cfg_din252,
   output        cfg_din253,
   output        cfg_din254,
   output        cfg_din255,
   output        cfg_din256,
   output        cfg_din257,
   output        cfg_din258,
   output        cfg_din259,
   output        cfg_din260,
   output        cfg_din261,
   output        cfg_din262,
   output        cfg_din263,
   output        cfg_din264,
   output        cfg_din265,
   output        cfg_din266,
   output        cfg_din267,
   output        cfg_din268,
   output        cfg_din269,
   output        cfg_din270,
   output        cfg_din271,
   output        cfg_din272,
   output        cfg_din273,
   output        cfg_din274,
   output        cfg_din275,
   output        cfg_din276,
   output        cfg_din277,
   output        cfg_din278,
   output        cfg_din279,
   output        cfg_din280,
   output        cfg_din281,
   output        cfg_din282,
   output        cfg_din283,
   output        cfg_din284,
   output        cfg_din285,
   output        cfg_din286,
   output        cfg_din287,
   output        cfg_din288,
   output        cfg_din289,
   output        cfg_din290,
   output        cfg_din291,
   output        cfg_din292,
   output        cfg_din293,
   output        cfg_din294,
   output        cfg_din295,
   output        cfg_din296,
   output        cfg_din297,
   output        cfg_din298,
   output        cfg_din299,
   output        cfg_din300,
   output        cfg_din301,
   output        cfg_din302,
   output        cfg_din303,
   output        cfg_din304,
   output        cfg_din305,
   output        cfg_din306,
   output        cfg_din307,
   output        cfg_din308,
   output        cfg_din309,
   output        cfg_din310,
   output        cfg_din311,
   output        cfg_din312,
   output        cfg_din313,
   output        cfg_din314,
   output        cfg_din315,
   output        cfg_din316,
   output        cfg_din317,
   output        cfg_din318,
   output        cfg_din319,
   output        cfg_din320,
   output        cfg_din321,
   output        cfg_din322,
   output        cfg_din323,
   output        cfg_din324,
   output        cfg_din325,
   output        cfg_din326,
   output        cfg_din327,
   output        cfg_din328,
   output        cfg_din329,
   output        cfg_din330,
   output        cfg_din331,
   output        cfg_din332,
   output        cfg_din333,
   output        cfg_din334,
   output        cfg_din335,
   output        cfg_din336,
   output        cfg_din337,
   output        cfg_din338,
   output        cfg_din339,
   output        cfg_din340,
   output        cfg_din341,
   output        cfg_din342,
   output        cfg_din343,
   output        cfg_din344,
   output        cfg_din345,
   output        cfg_din346,
   output        cfg_din347,
   output        cfg_din348,
   output        cfg_din349,
   output        cfg_din350,
   output        cfg_din351,
   output        cfg_din352,
   output        cfg_din353,
   output        cfg_din354,
   output        cfg_din355,
   output        cfg_din356,
   output        cfg_din357,
   output        cfg_din358,
   output        cfg_din359,
   output        cfg_din360,
   output        cfg_din361,
   output        cfg_din362,
   output        cfg_din363,
   output        cfg_din364,
   output        cfg_din365,
   output        cfg_din366,
   output        cfg_din367,
   output        cfg_din368,
   output        cfg_din369,
   output        cfg_din370,
   output        cfg_din371,
   output        cfg_din372,
   output        cfg_din373,
   output        cfg_din374,
   output        cfg_din375,
   output        cfg_din376,
   output        cfg_din377,
   output        cfg_din378,
   output        cfg_din379,
   output        cfg_din380,
   output        cfg_din381,
   output        cfg_din382,
   output        cfg_din383,
   output        cfg_din384,
   output        cfg_din385,
   output        cfg_din386,
   output        cfg_din387,
   output        cfg_din388,
   output        cfg_din389,
   output        cfg_din390,
   output        cfg_din391,
   output        cfg_din392,
   output        cfg_din393,
   output        cfg_din394,
   output        cfg_din395,
   output        cfg_din396,
   output        cfg_din397,
   output        cfg_din398,
   output        cfg_din399,
   output        cfg_din400,
   output        cfg_din401,
   output        cfg_din402,
   output        cfg_din403,
   output        cfg_din404,
   output        cfg_din405,
   output        cfg_din406,
   output        cfg_din407,
   output        cfg_din408,
   output        cfg_din409,
   output        cfg_din410,
   output        cfg_din411,
   output        cfg_din412,
   output        cfg_din413,
   output        cfg_din414,
   output        cfg_din415,
   output        cfg_din416,
   output        cfg_din417,
   output        cfg_din418,
   output        cfg_din419,
   output        cfg_din420,
   output        cfg_din421,
   output        cfg_din422,
   output        cfg_din423,
   output        cfg_din424,
   output        cfg_din425,
   output        cfg_din426,
   output        cfg_din427,
   output        cfg_din428,
   output        cfg_din429,
   output        cfg_din430,
   output        cfg_din431,
   output        cfg_din432,
   output        cfg_din433,
   output        cfg_din434,
   output        cfg_din435,
   output        cfg_din436,
   output        cfg_din437,
   output        cfg_din438,
   output        cfg_din439,
   output        cfg_din440,
   output        cfg_din441,
   output        cfg_din442,
   output        cfg_din443,
   output        cfg_din444,
   output        cfg_din445,
   output        cfg_din446,
   output        cfg_din447,
   output        cfg_din448,
   output        cfg_din449,
   output        cfg_din450,
   output        cfg_din451,
   output        cfg_din452,
   output        cfg_din453,
   output        cfg_din454,
   output        cfg_din455,
   output        cfg_din456,
   output        cfg_din457,
   output        cfg_din458,
   output        cfg_din459,
   output        cfg_din460,
   output        cfg_din461,
   output        cfg_din462,
   output        cfg_din463,
   output        cfg_din464,
   output        cfg_din465,
   output        cfg_din466,
   output        cfg_din467,
   output        cfg_din468,
   output        cfg_din469,
   output        cfg_din470,
   output        cfg_din471,
   output        cfg_din472,
   output        cfg_din473,
   output        cfg_din474,
   output        cfg_din475,
   output        cfg_din476,
   output        cfg_din477,
   output        cfg_din478,
   output        cfg_din479,
   output        cfg_din480,
   output        cfg_din481,
   output        cfg_din482,
   output        cfg_din483,
   output        cfg_din484,
   output        cfg_din485,
   output        cfg_din486,
   output        cfg_din487,
   output        cfg_din488,
   output        cfg_din489,
   output        cfg_din490,
   output        cfg_din491,
   output        cfg_din492,
   output        cfg_din493,
   output        cfg_din494,
   output        cfg_din495,
   output        cfg_din496,
   output        cfg_din497,
   output        cfg_din498,
   output        cfg_din499,
   output        cfg_din500,
   output        cfg_din501,
   output        cfg_din502,
   output        cfg_din503,
   output        cfg_din504,
   output        cfg_din505,
   output        cfg_din506,
   output        cfg_din507,
   output        cfg_din508,
   output        cfg_din509,
   output        cfg_din510,
   output        cfg_din511,
   output        cfg_din512,
   output        cfg_din513,
   output        cfg_din514,
   output        cfg_din515,
   output        cfg_din516,
   output        cfg_din517,
   output        cfg_din518,
   output        cfg_din519,
   output        cfg_din520,
   output        cfg_din521,
   output        cfg_din522,
   output        cfg_din523,
   output        cfg_din524,
   output        cfg_din525,
   output        cfg_din526,
   output        cfg_din527,
   output        cfg_din528,
   output        cfg_din529,
   output        cfg_din530,
   output        cfg_din531,
   output        cfg_din532,
   output        cfg_din533,
   output        cfg_din534,
   output        cfg_din535,
   output        cfg_din536,
   output        cfg_din537,
   output        cfg_din538,
   output        cfg_din539,
   output        cfg_din540,
   output        cfg_din541,
   output        cfg_din542,
   output        cfg_din543,
   output        cfg_din544,
   output        cfg_din545,
   output        cfg_din546,
   output        cfg_din547,
   output        cfg_din548,
   output        cfg_din549,
   output        cfg_din550,
   output        cfg_din551,
   output        cfg_din552,
   output        cfg_din553,
   output        cfg_din554,
   output        cfg_din555,
   output        cfg_din556,
   output        cfg_din557,
   output        cfg_din558,
   output        cfg_din559,
   output        cfg_din560,
   output        cfg_din561,
   output        cfg_din562,
   output        cfg_din563,
   output        cfg_din564,
   output        cfg_din565,
   output        cfg_din566,
   output        cfg_din567,
   output        cfg_din568,
   output        cfg_din569,
   output        cfg_din570,
   output        cfg_din571,
   output        cfg_din572,
   output        cfg_din573,
   output        cfg_din574,
   output        cfg_din575,
   output        cfg_din576,
   output        cfg_din577,
   output        cfg_din578,
   output        cfg_din579,
   output        cfg_din580,
   output        cfg_din581,
   output        cfg_din582,
   output        cfg_din583,
   output        cfg_din584,
   output        cfg_din585,
   output        cfg_din586,
   output        cfg_din587,
   output        cfg_din588,
   output        cfg_din589,
   output        cfg_din590,
   output        cfg_din591,
   output        cfg_din592,
   output        cfg_din593,
   output        cfg_din594,
   output        cfg_din595,
   output        cfg_din596,
   output        cfg_din597,
   output        cfg_din598,
   output        cfg_din599,
   output        cfg_din600,
   output        cfg_din601,
   output        cfg_din602,
   output        cfg_din603,
   output        cfg_din604,
   output        cfg_din605,
   output        cfg_din606,
   output        cfg_din607,
   output        cfg_din608,
   output        cfg_din609,
   output        cfg_din610,
   output        cfg_din611,
   output        cfg_din612,
   output        cfg_din613,
   output        cfg_din614,
   output        cfg_din615,
   output        cfg_din616,
   output        cfg_din617,
   output        cfg_din618,
   output        cfg_din619,
   output        cfg_din620,
   output        cfg_din621,
   output        cfg_din622,
   output        cfg_din623,
   output        cfg_din624,
   output        cfg_din625,
   output        cfg_din626,
   output        cfg_din627,
   output        cfg_din628,
   output        cfg_din629,
   output        cfg_din630,
   output        cfg_din631,
   output        cfg_din632,
   output        cfg_din633,
   output        cfg_din634,
   output        cfg_din635,
   output        cfg_din636,
   output        cfg_din637,
   output        cfg_din638,
   output        cfg_din639,
   output        cfg_din640,
   output        cfg_din641,
   output        cfg_din642,
   output        cfg_din643,
   output        cfg_din644,
   output        cfg_din645,
   output        cfg_din646,
   output        cfg_din647,
   output        cfg_din648,
   output        cfg_din649,
   output        cfg_din650,
   output        cfg_din651,
   output        cfg_din652,
   output        cfg_din653,
   output        cfg_din654,
   output        cfg_din655,
   output        cfg_din656,
   output        cfg_din657,
   output        cfg_din658,
   output        cfg_din659,
   output        cfg_din660,
   output        cfg_din661,
   output        cfg_din662,
   output        cfg_din663,
   output        cfg_din664,
   output        cfg_din665,
   output        cfg_din666,
   output        cfg_din667,
   output        cfg_din668,
   output        cfg_din669,
   output        cfg_din670,
   output        cfg_din671,
   output        cfg_din672,
   output        cfg_din673,
   output        cfg_din674,
   output        cfg_din675,
   output        cfg_din676,
   output        cfg_din677,
   output        cfg_din678,
   output        cfg_din679,
   output        cfg_din680,
   output        cfg_din681,
   output        cfg_din682,
   output        cfg_din683,
   output        cfg_din684,
   output        cfg_din685,
   output        cfg_din686,
   output        cfg_din687,
   output        cfg_din688,
   output        cfg_din689,
   output        cfg_din690,
   output        cfg_din691,
   output        cfg_din692,
   output        cfg_din693,
   output        cfg_din694,
   output        cfg_din695,
   output        cfg_din696,
   output        cfg_din697,
   output        cfg_din698,
   output        cfg_din699,
   output        cfg_din700,
   output        cfg_din701,
   output        cfg_din702,
   output        cfg_din703,
   output        cfg_din704,
   output        cfg_din705,
   output        cfg_din706,
   output        cfg_din707,
   output        cfg_din708,
   output        cfg_din709,
   output        cfg_din710,
   output        cfg_din711,
   output        cfg_din712,
   output        cfg_din713,
   output        cfg_din714,
   output        cfg_din715,
   output        cfg_din716,
   output        cfg_din717,
   output        cfg_din718,
   output        cfg_din719,
   output        cfg_din720,
   output        cfg_din721,
   output        cfg_din722,
   output        cfg_din723,
   output        cfg_din724,
   output        cfg_din725,
   output        cfg_din726,
   output        cfg_din727,
   output        cfg_din728,
   output        cfg_din729,
   output        cfg_din730,
   output        cfg_din731,
   output        cfg_din732,
   output        cfg_din733,
   output        cfg_din734,
   output        cfg_din735,
   output        cfg_din736,
   output        cfg_din737,
   output        cfg_din738,
   output        cfg_din739,
   output        cfg_din740,
   output        cfg_din741,
   output        cfg_din742,
   output        cfg_din743,
   output        cfg_din744,
   output        cfg_din745,
   output        cfg_din746,
   output        cfg_din747,
   output        cfg_din748,
   output        cfg_din749,
   output        cfg_din750,
   output        cfg_din751,
   output        cfg_din752,
   output        cfg_din753,
   output        cfg_din754,
   output        cfg_din755,
   output        cfg_din756,
   output        cfg_din757,
   output        cfg_din758,
   output        cfg_din759,
   output        cfg_din760,
   output        cfg_din761,
   output        cfg_din762,
   output        cfg_din763,
   output        cfg_din764,
   output        cfg_din765,
   output        cfg_din766,
   output        cfg_din767,
   output        cfg_din768,
   output        cfg_din769,
   output        cfg_din770,
   output        cfg_din771,
   output        cfg_din772,
   output        cfg_din773,
   output        cfg_din774,
   output        cfg_din775,
   output        cfg_din776,
   output        cfg_din777,
   output        cfg_din778,
   output        cfg_din779,
   output        cfg_din780,
   output        cfg_din781,
   output        cfg_din782,
   output        cfg_din783,
   output        cfg_din784,
   output        cfg_din785,
   output        cfg_din786,
   output        cfg_din787,
   output        cfg_din788,
   output        cfg_din789,
   output        cfg_din790,
   output        cfg_din791,
   output        cfg_din792,
   output        cfg_din793,
   output        cfg_din794,
   output        cfg_din795,
   output        cfg_din796,
   output        cfg_din797,
   output        cfg_din798,
   output        cfg_din799,
   output        cfg_din800,
   output        cfg_din801,
   output        cfg_din802,
   output        cfg_din803,
   output        cfg_din804,
   output        cfg_din805,
   output        cfg_din806,
   output        cfg_din807,
   output        cfg_din808,
   output        cfg_din809,
   output        cfg_din810,
   output        cfg_din811,
   output        cfg_din812,
   output        cfg_din813,
   output        cfg_din814,
   output        cfg_din815,
   output        cfg_din816,
   output        cfg_din817,
   output        cfg_din818,
   output        cfg_din819,
   output        cfg_din820,
   output        cfg_din821,
   output        cfg_din822,
   output        cfg_din823,
   output        cfg_din824,
   output        cfg_din825,
   output        cfg_din826,
   output        cfg_din827,
   output        cfg_din828,
   output        cfg_din829,
   output        cfg_din830,
   output        cfg_din831,
   output        cfg_din832,
   output        cfg_din833,
   output        cfg_din834,
   output        cfg_din835,
   output        cfg_din836,
   output        cfg_din837,
   output        cfg_din838,
   output        cfg_din839,
   output        cfg_din840,
   output        cfg_din841,
   output        cfg_din842,
   output        cfg_din843,
   output        cfg_din844,
   output        cfg_din845,
   output        cfg_din846,
   output        cfg_din847,
   output        cfg_din848,
   output        cfg_din849,
   output        cfg_din850,
   output        cfg_din851,
   output        cfg_din852,
   output        cfg_din853,
   output        cfg_din854,
   output        cfg_din855,
   output        cfg_din856,
   output        cfg_din857,
   output        cfg_din858,
   output        cfg_din859,
   output        cfg_din860,
   output        cfg_din861,
   output        cfg_din862,
   output        cfg_din863,
   output        cfg_din864,
   output        cfg_din865,
   output        cfg_din866,
   output        cfg_din867,
   output        cfg_din868,
   output        cfg_din869,
   output        cfg_din870,
   output        cfg_din871,
   output        cfg_din872,
   output        cfg_din873,
   output        cfg_din874,
   output        cfg_din875,
   output        cfg_din876,
   output        cfg_din877,
   output        cfg_din878,
   output        cfg_din879,
   output        cfg_din880,
   output        cfg_din881,
   output        cfg_din882,
   output        cfg_din883,
   output        cfg_din884,
   output        cfg_din885,
   output        cfg_din886,
   output        cfg_din887,
   output        cfg_din888,
   output        cfg_din889,
   output        cfg_din890,
   output        cfg_din891,
   output        cfg_din892,
   output        cfg_din893,
   output        cfg_din894,
   output        cfg_din895,
   output        cfg_din896,
   output        cfg_din897,
   output        cfg_din898,
   output        cfg_din899,
   output        cfg_din900,
   output        cfg_din901,
   output        cfg_din902,
   output        cfg_din903,
   output        cfg_din904,
   output        cfg_din905,
   output        cfg_din906,
   output        cfg_din907,
   output        cfg_din908,
   output        cfg_din909,
   output        cfg_din910,
   output        cfg_din911,
   output        cfg_din912,
   output        cfg_din913,
   output        cfg_din914,
   output        cfg_din915,
   output        cfg_din916,
   output        cfg_din917,
   output        cfg_din918,
   output        cfg_din919,
   output        cfg_din920,
   output        cfg_din921,
   output        cfg_din922,
   output        cfg_din923,
   output        cfg_din924,
   output        cfg_din925,
   output        cfg_din926,
   output        cfg_din927,
   output        cfg_din928,
   output        cfg_din929,
   output        cfg_din930,
   output        cfg_din931,
   output        cfg_din932,
   output        cfg_din933,
   output        cfg_din934,
   output        cfg_din935,
   output        cfg_din936,
   output        cfg_din937,
   output        cfg_din938,
   output        cfg_din939,
   output        cfg_din940,
   output        cfg_din941,
   output        cfg_din942,
   output        cfg_din943,
   output        cfg_din944,
   output        cfg_din945,
   output        cfg_din946,
   output        cfg_din947,
   output        cfg_din948,
   output        cfg_din949,
   output        cfg_din950,
   output        cfg_din951,
   output        cfg_din952,
   output        cfg_din953,
   output        cfg_din954,
   output        cfg_din955,
   output        cfg_din956,
   output        cfg_din957,
   output        cfg_din958,
   output        cfg_din959,
   output        cfg_din960,
   output        cfg_din961,
   output        cfg_din962,
   output        cfg_din963,
   output        cfg_din964,
   output        cfg_din965,
   output        cfg_din966,
   output        cfg_din967,
   output        cfg_din968,
   output        cfg_din969,
   output        cfg_din970,
   output        cfg_din971,
   output        cfg_din972,
   output        cfg_din973,
   output        cfg_din974,
   output        cfg_din975,
   output        cfg_din976,
   output        cfg_din977,
   output        cfg_din978,
   output        cfg_din979,
   output        cfg_din980,
   output        cfg_din981,
   output        cfg_din982,
   output        cfg_din983,
   output        cfg_din984,
   output        cfg_din985,
   output        cfg_din986,
   output        cfg_din987,
   output        cfg_din988,
   output        cfg_din989,
   output        cfg_din990,
   output        cfg_din991,
   output        cfg_din992,
   output        cfg_din993,
   output        cfg_din994,
   output        cfg_din995,
   output        cfg_din996,
   output        cfg_din997,
   output        cfg_din998,
   output        cfg_din999,
   output        cfg_din1000,
   output        cfg_din1001,
   output        cfg_din1002,
   output        cfg_din1003,
   output        cfg_din1004,
   output        cfg_din1005,
   output        cfg_din1006,
   output        cfg_din1007,
   output        cfg_din1008,
   output        cfg_din1009,
   output        cfg_din1010,
   output        cfg_din1011,
   output        cfg_din1012,
   output        cfg_din1013,
   output        cfg_din1014,
   output        cfg_din1015,
   output        cfg_din1016,
   output        cfg_din1017,
   output        cfg_din1018,
   output        cfg_din1019,
   output        cfg_din1020,
   output        cfg_din1021,
   output        cfg_din1022,
   output        cfg_din1023,
   output        cfg_din1024,
   output        cfg_din1025,
   output        cfg_din1026,
   output        cfg_din1027,
   output        cfg_din1028,
   output        cfg_din1029,
   output        cfg_din1030,
   output        cfg_din1031,
   output        cfg_din1032,
   output        cfg_din1033,
   output        cfg_din1034,
   output        cfg_din1035,
   output        cfg_din1036,
   output        cfg_din1037,
   output        cfg_din1038,
   output        cfg_din1039,
   output        cfg_din1040,
   output        cfg_din1041,
   output        cfg_din1042,
   output        cfg_din1043,
   output        cfg_din1044,
   output        cfg_din1045,
   output        cfg_din1046,
   output        cfg_din1047,
   output        cfg_din1048,
   output        cfg_din1049,
   output        cfg_din1050,
   output        cfg_din1051,
   output        cfg_din1052,
   output        cfg_din1053,
   output        cfg_din1054,
   output        cfg_din1055,
   output        cfg_din1056,
   output        cfg_din1057,
   output        cfg_din1058,
   output        cfg_din1059,
   output        cfg_din1060,
   output        cfg_din1061,
   output        cfg_din1062,
   output        cfg_din1063,
   output        cfg_din1064,
   output        cfg_din1065,
   output        cfg_din1066,
   output        cfg_din1067,
   output        cfg_din1068,
   output        cfg_din1069,
   output        cfg_din1070,
   output        cfg_din1071,
   output        cfg_din1072,
   output        cfg_din1073,
   output        cfg_din1074,
   output        cfg_din1075,
   output        cfg_din1076,
   output        cfg_din1077,
   output        cfg_din1078,
   output        cfg_din1079,
   output        cfg_din1080,
   output        cfg_din1081,
   output        cfg_din1082,
   output        cfg_din1083,
   output        cfg_din1084,
   output        cfg_din1085,
   output        cfg_din1086,
   output        cfg_din1087,
   output        cfg_din1088,
   output        cfg_din1089,
   output        cfg_din1090,
   output        cfg_din1091,
   output        cfg_din1092,
   output        cfg_din1093,
   output        cfg_din1094,
   output        cfg_din1095,
   output        cfg_din1096,
   output        cfg_din1097,
   output        cfg_din1098,
   output        cfg_din1099,
   output        cfg_din1100,
   output        cfg_din1101,
   output        cfg_din1102,
   output        cfg_din1103,
   output        cfg_din1104,
   output        cfg_din1105,
   output        cfg_din1106,
   output        cfg_din1107,
   output        cfg_din1108,
   output        cfg_din1109,
   output        cfg_din1110,
   output        cfg_din1111,
   output        cfg_din1112,
   output        cfg_din1113,
   output        cfg_din1114,
   output        cfg_din1115,
   output        cfg_din1116,
   output        cfg_din1117,
   output        cfg_din1118,
   output        cfg_din1119,
   output        cfg_din1120,
   output        cfg_din1121,
   output        cfg_din1122,
   output        cfg_din1123,
   output        cfg_din1124,
   output        cfg_din1125,
   output        cfg_din1126,
   output        cfg_din1127,
   output        cfg_din1128,
   output        cfg_din1129,
   output        cfg_din1130,
   output        cfg_din1131,
   output        cfg_din1132,
   output        cfg_din1133,
   output        cfg_din1134,
   output        cfg_din1135,
   output        cfg_din1136,
   output        cfg_din1137,
   output        cfg_din1138,
   output        cfg_din1139,
   output        cfg_din1140,
   output        cfg_din1141,
   output        cfg_din1142,
   output        cfg_din1143,
   output        cfg_din1144,
   output        cfg_din1145,
   output        cfg_din1146,
   output        cfg_din1147,
   output        cfg_din1148,
   output        cfg_din1149,
   output        cfg_din1150,
   output        cfg_din1151,
   output        cfg_din1152,
   output        cfg_din1153,
   output        cfg_din1154,
   output        cfg_din1155,
   output        cfg_din1156,
   output        cfg_din1157,
   output        cfg_din1158,
   output        cfg_din1159,
   output        cfg_din1160,
   output        cfg_din1161,
   output        cfg_din1162,
   output        cfg_din1163,
   output        cfg_din1164,
   output        cfg_din1165,
   output        cfg_din1166,
   output        cfg_din1167,
   output        cfg_din1168,
   output        cfg_din1169,
   output        cfg_din1170,
   output        cfg_din1171,
   output        cfg_din1172,
   output        cfg_din1173,
   output        cfg_din1174,
   output        cfg_din1175,
   output        cfg_din1176,
   output        cfg_din1177,
   output        cfg_din1178,
   output        cfg_din1179,
   output        cfg_din1180,
   output        cfg_din1181,
   output        cfg_din1182,
   output        cfg_din1183,
   output        cfg_din1184,
   output        cfg_din1185,
   output        cfg_din1186,
   output        cfg_din1187,
   output        cfg_din1188,
   output        cfg_din1189,
   output        cfg_din1190,
   output        cfg_din1191,
   output        cfg_din1192,
   output        cfg_din1193,
   output        cfg_din1194,
   output        cfg_din1195,
   output        cfg_din1196,
   output        cfg_din1197,
   output        cfg_din1198,
   output        cfg_din1199,
   output        cfg_din1200,
   output        cfg_din1201,
   output        cfg_din1202,
   output        cfg_din1203,
   output        cfg_din1204,
   output        cfg_din1205,
   output        cfg_din1206,
   output        cfg_din1207,
   output        cfg_din1208,
   output        cfg_din1209,
   output        cfg_din1210,
   output        cfg_din1211,
   output        cfg_din1212,
   output        cfg_din1213,
   output        cfg_din1214,
   output        cfg_din1215,
   output        cfg_din1216,
   output        cfg_din1217,
   output        cfg_din1218,
   output        cfg_din1219,
   output        cfg_din1220,
   output        cfg_din1221,
   output        cfg_din1222,
   output        cfg_din1223,
   output        cfg_din1224,
   output        cfg_din1225,
   output        cfg_din1226,
   output        cfg_din1227,
   output        cfg_din1228,
   output        cfg_din1229,
   output        cfg_din1230,
   output        cfg_din1231,
   output        cfg_din1232,
   output        cfg_din1233,
   output        cfg_din1234,
   output        cfg_din1235,
   output        cfg_din1236,
   output        cfg_din1237,
   output        cfg_din1238,
   output        cfg_din1239,
   output        cfg_din1240,
   output        cfg_din1241,
   output        cfg_din1242,
   output        cfg_din1243,
   output        cfg_din1244,
   output        cfg_din1245,
   output        cfg_din1246,
   output        cfg_din1247,
   output        cfg_din1248,
   output        cfg_din1249,
   output        cfg_din1250,
   output        cfg_din1251,
   output        cfg_din1252,
   output        cfg_din1253,
   output        cfg_din1254,
   output        cfg_din1255,
   output        cfg_din1256,
   output        cfg_din1257,
   output        cfg_din1258,
   output        cfg_din1259,
   output        cfg_din1260,
   output        cfg_din1261,
   output        cfg_din1262,
   output        cfg_din1263,
   output        cfg_din1264,
   output        cfg_din1265,
   output        cfg_din1266,
   output        cfg_din1267,
   output        cfg_din1268,
   output        cfg_din1269,
   output        cfg_din1270,
   output        cfg_din1271,
   output        cfg_din1272,
   output        cfg_din1273,
   output        cfg_din1274,
   output        cfg_din1275,
   output        cfg_din1276,
   output        cfg_din1277,
   output        cfg_din1278,
   output        cfg_din1279,
   output        cfg_din1280,
   output        cfg_din1281,
   output        cfg_din1282,
   output        cfg_din1283,
   output        cfg_din1284,
   output        cfg_din1285,
   output        cfg_din1286,
   output        cfg_din1287,
   output        cfg_din1288,
   output        cfg_din1289,
   output        cfg_din1290,
   output        cfg_din1291,
   output        cfg_din1292,
   output        cfg_din1293,
   output        cfg_din1294,
   output        cfg_din1295,
   output        cfg_din1296,
   output        cfg_din1297,
   output        cfg_din1298,
   output        cfg_din1299,
   output        cfg_din1300,
   output        cfg_din1301,
   output        cfg_din1302,
   output        cfg_din1303,
   output        cfg_din1304,
   output        cfg_din1305,
   output        cfg_din1306,
   output        cfg_din1307,
   output        cfg_din1308,
   output        cfg_din1309,
   output        cfg_din1310,
   output        cfg_din1311,
   output        cfg_din1312,
   output        cfg_din1313,
   output        cfg_din1314,
   output        cfg_din1315,
   output        cfg_din1316,
   output        cfg_din1317,
   output        cfg_din1318,
   output        cfg_din1319,
   output        cfg_din1320,
   output        cfg_din1321,
   output        cfg_din1322,
   output        cfg_din1323,
   output        cfg_din1324,
   output        cfg_din1325,
   output        cfg_din1326,
   output        cfg_din1327,
   output        cfg_din1328,
   output        cfg_din1329,
   output        cfg_din1330,
   output        cfg_din1331,
   output        cfg_din1332,
   output        cfg_din1333,
   output        cfg_din1334,
   output        cfg_din1335,
   output        cfg_din1336,
   output        cfg_din1337,
   output        cfg_din1338,
   output        cfg_din1339,
   output        cfg_din1340,
   output        cfg_din1341,
   output        cfg_din1342,
   output        cfg_din1343,
   output        cfg_din1344,
   output        cfg_din1345,
   output        cfg_din1346,
   output        cfg_din1347,
   output        cfg_din1348,
   output        cfg_din1349,
   output        cfg_din1350,
   output        cfg_din1351,
   output        cfg_din1352,
   output        cfg_din1353,
   output        cfg_din1354,
   output        cfg_din1355,
   output        cfg_din1356,
   output        cfg_din1357,
   output        cfg_din1358,
   output        cfg_din1359,
   output        cfg_din1360,
   output        cfg_din1361,
   output        cfg_din1362,
   output        cfg_din1363,
   output        cfg_din1364,
   output        cfg_din1365,
   output        cfg_din1366,
   output        cfg_din1367,
   output        cfg_din1368,
   output        cfg_din1369,
   output        cfg_din1370,
   output        cfg_din1371,
   output        cfg_din1372,
   output        cfg_din1373,
   output        cfg_din1374,
   output        cfg_din1375,
   output        cfg_din1376,
   output        cfg_din1377,
   output        cfg_din1378,
   output        cfg_din1379,
   output        cfg_din1380,
   output        cfg_din1381,
   output        cfg_din1382,
   output        cfg_din1383,
   output        cfg_din1384,
   output        cfg_din1385,
   output        cfg_din1386,
   output        cfg_din1387,
   output        cfg_din1388,
   output        cfg_din1389,
   output        cfg_din1390,
   output        cfg_din1391,
   output        cfg_din1392,
   output        cfg_din1393,
   output        cfg_din1394,
   output        cfg_din1395,
   output        cfg_din1396,
   output        cfg_din1397,
   output        cfg_din1398,
   output        cfg_din1399,
   output        cfg_din1400,
   output        cfg_din1401,
   output        cfg_din1402,
   output        cfg_din1403,
   output        cfg_din1404,
   output        cfg_din1405,
   output        cfg_din1406,
   output        cfg_din1407,
   output        cfg_din1408,
   output        cfg_din1409,
   output        cfg_din1410,
   output        cfg_din1411,
   output        cfg_din1412,
   output        cfg_din1413,
   output        cfg_din1414,
   output        cfg_din1415,
   output        cfg_din1416,
   output        cfg_din1417,
   output        cfg_din1418,
   output        cfg_din1419,
   output        cfg_din1420,
   output        cfg_din1421,
   output        cfg_din1422,
   output        cfg_din1423,
   output        cfg_din1424,
   output        cfg_din1425,
   output        cfg_din1426,
   output        cfg_din1427,
   output        cfg_din1428,
   output        cfg_din1429,
   output        cfg_din1430,
   output        cfg_din1431,
   output        cfg_din1432,
   output        cfg_din1433,
   output        cfg_din1434,
   output        cfg_din1435,
   output        cfg_din1436,
   output        cfg_din1437,
   output        cfg_din1438,
   output        cfg_din1439,
   output        cfg_din1440,
   output        cfg_din1441,
   output        cfg_din1442,
   output        cfg_din1443,
   output        cfg_din1444,
   output        cfg_din1445,
   output        cfg_din1446,
   output        cfg_din1447,
   output        cfg_din1448,
   output        cfg_din1449,
   output        cfg_din1450,
   output        cfg_din1451,
   output        cfg_din1452,
   output        cfg_din1453,
   output        cfg_din1454,
   output        cfg_din1455,
   output        cfg_din1456,
   output        cfg_din1457,
   output        cfg_din1458,
   output        cfg_din1459,
   output        cfg_din1460,
   output        cfg_din1461,
   output        cfg_din1462,
   output        cfg_din1463,
   output        cfg_din1464,
   output        cfg_din1465,
   output        cfg_din1466,
   output        cfg_din1467,
   output        cfg_din1468,
   output        cfg_din1469,
   output        cfg_din1470,
   output        cfg_din1471,
   output        cfg_din1472,
   output        cfg_din1473,
   output        cfg_din1474,
   output        cfg_din1475,
   output        cfg_din1476,
   output        cfg_din1477,
   output        cfg_din1478,
   output        cfg_din1479,
   output        cfg_din1480,
   output        cfg_din1481,
   output        cfg_din1482,
   output        cfg_din1483,
   output        cfg_din1484,
   output        cfg_din1485,
   output        cfg_din1486,
   output        cfg_din1487,
   output        cfg_din1488,
   output        cfg_din1489,
   output        cfg_din1490,
   output        cfg_din1491,
   output        cfg_din1492,
   output        cfg_din1493,
   output        cfg_din1494,
   output        cfg_din1495,
   output        cfg_din1496,
   output        cfg_din1497,
   output        cfg_din1498,
   output        cfg_din1499,
   output        cfg_din1500,
   output        cfg_din1501,
   output        cfg_din1502,
   output        cfg_din1503,
   output        cfg_din1504,
   output        cfg_din1505,
   output        cfg_din1506,
   output        cfg_din1507,
   output        cfg_din1508,
   output        cfg_din1509,
   output        cfg_din1510,
   output        cfg_din1511,
   output        cfg_din1512,
   output        cfg_din1513,
   output        cfg_din1514,
   output        cfg_din1515,
   output        cfg_din1516,
   output        cfg_din1517,
   output        cfg_din1518,
   output        cfg_din1519,
   output        cfg_din1520,
   output        cfg_din1521,
   output        cfg_din1522,
   output        cfg_din1523,
   output        cfg_din1524,
   output        cfg_din1525,
   output        cfg_din1526,
   output        cfg_din1527,
   output        cfg_din1528,
   output        cfg_din1529,
   output        cfg_din1530,
   output        cfg_din1531,
   output        cfg_din1532,
   output        cfg_din1533,
   output        cfg_din1534,
   output        cfg_din1535,
   output        cfg_din1536,
   output        cfg_din1537,
   output        cfg_din1538,
   output        cfg_din1539,
   output        cfg_din1540,
   output        cfg_din1541,
   output        cfg_din1542,
   output        cfg_din1543,
   output        cfg_din1544,
   output        cfg_din1545,
   output        cfg_din1546,
   output        cfg_din1547,
   output        cfg_din1548,
   output        cfg_din1549,
   output        cfg_din1550,
   output        cfg_din1551,
   output        cfg_din1552,
   output        cfg_din1553,
   output        cfg_din1554,
   output        cfg_din1555,
   output        cfg_din1556,
   output        cfg_din1557,
   output        cfg_din1558,
   output        cfg_din1559,
   output        cfg_din1560,
   output        cfg_din1561,
   output        cfg_din1562,
   output        cfg_din1563,
   output        cfg_din1564,
   output        cfg_din1565,
   output        cfg_din1566,
   output        cfg_din1567,
   output        cfg_din1568,
   output        cfg_din1569,
   output        cfg_din1570,
   output        cfg_din1571,
   output        cfg_din1572,
   output        cfg_din1573,
   output        cfg_din1574,
   output        cfg_din1575,
   output        cfg_din1576,
   output        cfg_din1577,
   output        cfg_din1578,
   output        cfg_din1579,
   output        cfg_din1580,
   output        cfg_din1581,
   output        cfg_din1582,
   output        cfg_din1583,
   output        cfg_din1584,
   output        cfg_din1585,
   output        cfg_din1586,
   output        cfg_din1587,
   output        cfg_din1588,
   output        cfg_din1589,
   output        cfg_din1590,
   output        cfg_din1591,
   output        cfg_din1592,
   output        cfg_din1593,
   output        cfg_din1594,
   output        cfg_din1595,
   output        cfg_din1596,
   output        cfg_din1597,
   output        cfg_din1598,
   output        cfg_din1599,
   output        cfg_din1600,
   output        cfg_din1601,
   output        cfg_din1602,
   output        cfg_din1603,
   output        cfg_din1604,
   output        cfg_din1605,
   output        cfg_din1606,
   output        cfg_din1607,
   output        cfg_din1608,
   output        cfg_din1609,
   output        cfg_din1610,
   output        cfg_din1611,
   output        cfg_din1612,
   output        cfg_din1613,
   output        cfg_din1614,
   output        cfg_din1615,
   output        cfg_din1616,
   output        cfg_din1617,
   output        cfg_din1618,
   output        cfg_din1619,
   output        cfg_din1620,
   output        cfg_din1621,
   output        cfg_din1622,
   output        cfg_din1623,
   output        cfg_din1624,
   output        cfg_din1625,
   output        cfg_din1626,
   output        cfg_din1627,
   output        cfg_din1628,
   output        cfg_din1629,
   output        cfg_din1630,
   output        cfg_din1631,
   output        cfg_din1632,
   output        cfg_din1633,
   output        cfg_din1634,
   output        cfg_din1635,
   output        cfg_din1636,
   output        cfg_din1637,
   output        cfg_din1638,
   output        cfg_din1639,
   output        cfg_din1640,
   output        cfg_din1641,
   output        cfg_din1642,
   output        cfg_din1643,
   output        cfg_din1644,
   output        cfg_din1645,
   output        cfg_din1646,
   output        cfg_din1647,
   output        cfg_din1648,
   output        cfg_din1649,
   output        cfg_din1650,
   output        cfg_din1651,
   output        cfg_din1652,
   output        cfg_din1653,
   output        cfg_din1654,
   output        cfg_din1655,
   output        cfg_din1656,
   output        cfg_din1657,
   output        cfg_din1658,
   output        cfg_din1659,
   output        cfg_din1660,
   output        cfg_din1661,
   output        cfg_din1662,
   output        cfg_din1663,
   output        cfg_din1664,
   output        cfg_din1665,
   output        cfg_din1666,
   output        cfg_din1667,
   output        cfg_din1668,
   output        cfg_din1669,
   output        cfg_din1670,
   output        cfg_din1671,
   output        cfg_din1672,
   output        cfg_din1673,
   output        cfg_din1674,
   output        cfg_din1675,
   output        cfg_din1676,
   output        cfg_din1677,
   output        cfg_din1678,
   output        cfg_din1679,
   output        cfg_din1680,
   output        cfg_din1681,
   output        cfg_din1682,
   output        cfg_din1683,
   output        cfg_din1684,
   output        cfg_din1685,
   output        cfg_din1686,
   output        cfg_din1687,
   output        cfg_din1688,
   output        cfg_din1689,
   output        cfg_din1690,
   output        cfg_din1691,
   output        cfg_din1692,
   output        cfg_din1693,
   output        cfg_din1694,
   output        cfg_din1695,
   output        cfg_din1696,
   output        cfg_din1697,
   output        cfg_din1698,
   output        cfg_din1699,
   output        cfg_din1700,
   output        cfg_din1701,
   output        cfg_din1702,
   output        cfg_din1703,
   output        cfg_din1704,
   output        cfg_din1705,
   output        cfg_din1706,
   output        cfg_din1707,
   output        cfg_din1708,
   output        cfg_din1709,
   output        cfg_din1710,
   output        cfg_din1711,
   output        cfg_din1712,
   output        cfg_din1713,
   output        cfg_din1714,
   output        cfg_din1715,
   output        cfg_din1716,
   output        cfg_din1717,
   output        cfg_din1718,
   output        cfg_din1719,
   output        cfg_din1720,
   output        cfg_din1721,
   output        cfg_din1722,
   output        cfg_din1723,
   output        cfg_din1724,
   output        cfg_din1725,
   output        cfg_din1726,
   output        cfg_din1727,
   output        cfg_din1728,
   output        cfg_din1729,
   output        cfg_din1730,
   output        cfg_din1731,
   output        cfg_din1732,
   output        cfg_din1733,
   output        cfg_din1734,
   output        cfg_din1735,
   output        cfg_din1736,
   output        cfg_din1737,
   output        cfg_din1738,
   output        cfg_din1739,
   output        cfg_din1740,
   output        cfg_din1741,
   output        cfg_din1742,
   output        cfg_din1743,
   output        cfg_din1744,
   output        cfg_din1745,
   output        cfg_din1746,
   output        cfg_din1747,
   output        cfg_din1748,
   output        cfg_din1749,
   output        cfg_din1750,
   output        cfg_din1751,
   output        cfg_din1752,
   output        cfg_din1753,
   output        cfg_din1754,
   output        cfg_din1755,
   output        cfg_din1756,
   output        cfg_din1757,
   output        cfg_din1758,
   output        cfg_din1759,
   output        cfg_din1760,
   output        cfg_din1761,
   output        cfg_din1762,
   output        cfg_din1763,
   output        cfg_din1764,
   output        cfg_din1765,
   output        cfg_din1766,
   output        cfg_din1767,
   output        cfg_din1768,
   output        cfg_din1769,
   output        cfg_din1770,
   output        cfg_din1771,
   output        cfg_din1772,
   output        cfg_din1773,
   output        cfg_din1774,
   output        cfg_din1775,
   output        cfg_din1776,
   output        cfg_din1777,
   output        cfg_din1778,
   output        cfg_din1779,
   output        cfg_din1780,
   output        cfg_din1781,
   output        cfg_din1782,
   output        cfg_din1783,
   output        cfg_din1784,
   output        cfg_din1785,
   output        cfg_din1786,
   output        cfg_din1787,
   output        cfg_din1788,
   output        cfg_din1789,
   output        cfg_din1790,
   output        cfg_din1791,
   output        cfg_din1792,
   output        cfg_din1793,
   output        cfg_din1794,
   output        cfg_din1795,
   output        cfg_din1796,
   output        cfg_din1797,
   output        cfg_din1798,
   output        cfg_din1799,
   output        cfg_din1800,
   output        cfg_din1801,
   output        cfg_din1802,
   output        cfg_din1803,
   output        cfg_din1804,
   output        cfg_din1805,
   output        cfg_din1806,
   output        cfg_din1807,
   output        cfg_din1808,
   output        cfg_din1809,
   output        cfg_din1810,
   output        cfg_din1811,
   output        cfg_din1812,
   output        cfg_din1813,
   output        cfg_din1814,
   output        cfg_din1815,
   output        cfg_din1816,
   output        cfg_din1817,
   output        cfg_din1818,
   output        cfg_din1819,
   output        cfg_din1820,
   output        cfg_din1821,
   output        cfg_din1822,
   output        cfg_din1823,
   output        cfg_din1824,
   output        cfg_din1825,
   output        cfg_din1826,
   output        cfg_din1827,
   output        cfg_din1828,
   output        cfg_din1829,
   output        cfg_din1830,
   output        cfg_din1831,
   output        cfg_din1832,
   output        cfg_din1833,
   output        cfg_din1834,
   output        cfg_din1835,
   output        cfg_din1836,
   output        cfg_din1837,
   output        cfg_din1838,
   output        cfg_din1839,
   output        cfg_din1840,
   output        cfg_din1841,
   output        cfg_din1842,
   output        cfg_din1843,
   output        cfg_din1844,
   output        cfg_din1845,
   output        cfg_din1846,
   output        cfg_din1847,
   output        cfg_din1848,
   output        cfg_din1849,
   output        cfg_din1850,
   output        cfg_din1851,
   output        cfg_din1852,
   output        cfg_din1853,
   output        cfg_din1854,
   output        cfg_din1855,
   output        cfg_din1856,
   output        cfg_din1857,
   output        cfg_din1858,
   output        cfg_din1859,
   output        cfg_din1860,
   output        cfg_din1861,
   output        cfg_din1862,
   output        cfg_din1863,
   output        cfg_din1864,
   output        cfg_din1865,
   output        cfg_din1866,
   output        cfg_din1867,
   output        cfg_din1868,
   output        cfg_din1869,
   output        cfg_din1870,
   output        cfg_din1871,
   output        cfg_din1872,
   output        cfg_din1873,
   output        cfg_din1874,
   output        cfg_din1875,
   output        cfg_din1876,
   output        cfg_din1877,
   output        cfg_din1878,
   output        cfg_din1879,
   output        cfg_din1880,
   output        cfg_din1881,
   output        cfg_din1882,
   output        cfg_din1883,
   output        cfg_din1884,
   output        cfg_din1885,
   output        cfg_din1886,
   output        cfg_din1887,
   output        cfg_din1888,
   output        cfg_din1889,
   output        cfg_din1890,
   output        cfg_din1891,
   output        cfg_din1892,
   output        cfg_din1893,
   output        cfg_din1894,
   output        cfg_din1895,
   output        cfg_din1896,
   output        cfg_din1897,
   output        cfg_din1898,
   output        cfg_din1899,
   output        cfg_din1900,
   output        cfg_din1901,
   output        cfg_din1902,
   output        cfg_din1903,
   output        cfg_din1904,
   output        cfg_din1905,
   output        cfg_din1906,
   output        cfg_din1907,
   output        cfg_din1908,
   output        cfg_din1909,
   output        cfg_din1910,
   output        cfg_din1911,
   output        cfg_din1912,
   output        cfg_din1913,
   output        cfg_din1914,
   output        cfg_din1915,
   output        cfg_din1916,
   output        cfg_din1917,
   output        cfg_din1918,
   output        cfg_din1919,
   output        cfg_din1920,
   output        cfg_din1921,
   output        cfg_din1922,
   output        cfg_din1923,
   output        cfg_din1924,
   output        cfg_din1925,
   output        cfg_din1926,
   output        cfg_din1927,
   output        cfg_din1928,
   output        cfg_din1929,
   output        cfg_din1930,
   output        cfg_din1931,
   output        cfg_din1932,
   output        cfg_din1933,
   output        cfg_din1934,
   output        cfg_din1935,
   output        cfg_din1936,
   output        cfg_din1937,
   output        cfg_din1938,
   output        cfg_din1939,
   output        cfg_din1940,
   output        cfg_din1941,
   output        cfg_din1942,
   output        cfg_din1943,
   output        cfg_din1944,
   output        cfg_din1945,
   output        cfg_din1946,
   output        cfg_din1947,
   output        cfg_din1948,
   output        cfg_din1949,
   output        cfg_din1950,
   output        cfg_din1951,
   output        cfg_din1952,
   output        cfg_din1953,
   output        cfg_din1954,
   output        cfg_din1955,
   output        cfg_din1956,
   output        cfg_din1957,
   output        cfg_din1958,
   output        cfg_din1959,
   output        cfg_din1960,
   output        cfg_din1961,
   output        cfg_din1962,
   output        cfg_din1963,
   output        cfg_din1964,
   output        cfg_din1965,
   output        cfg_din1966,
   output        cfg_din1967,
   output        cfg_din1968,
   output        cfg_din1969,
   output        cfg_din1970,
   output        cfg_din1971,
   output        cfg_din1972,
   output        cfg_din1973,
   output        cfg_din1974,
   output        cfg_din1975,
   output        cfg_din1976,
   output        cfg_din1977,
   output        cfg_din1978,
   output        cfg_din1979,
   output        cfg_din1980,
   output        cfg_din1981,
   output        cfg_din1982,
   output        cfg_din1983,
   output        cfg_din1984,
   output        cfg_din1985,
   output        cfg_din1986,
   output        cfg_din1987,
   output        cfg_din1988,
   output        cfg_din1989,
   output        cfg_din1990,
   output        cfg_din1991,
   output        cfg_din1992,
   output        cfg_din1993,
   output        cfg_din1994,
   output        cfg_din1995,
   output        cfg_din1996,
   output        cfg_din1997,
   output        cfg_din1998,
   output        cfg_din1999,
   output        cfg_din2000,
   output        cfg_din2001,
   output        cfg_din2002,
   output        cfg_din2003,
   output        cfg_din2004,
   output        cfg_din2005,
   output        cfg_din2006,
   output        cfg_din2007,
   output        cfg_din2008,
   output        cfg_din2009,
   output        cfg_din2010,
   output        cfg_din2011,
   output        cfg_din2012,
   output        cfg_din2013,
   output        cfg_din2014,
   output        cfg_din2015,
   output        cfg_din2016,
   output        cfg_din2017,
   output        cfg_din2018,
   output        cfg_din2019,
   output        cfg_din2020,
   output        cfg_din2021,
   output        cfg_din2022,
   output        cfg_din2023,
   output        cfg_din2024,
   output        cfg_din2025,
   output        cfg_din2026,
   output        cfg_din2027,
   output        cfg_din2028,
   output        cfg_din2029,
   output        cfg_din2030,
   output        cfg_din2031,
   output        cfg_din2032,
   output        cfg_din2033,
   output        cfg_din2034,
   output        cfg_din2035,
   output        cfg_din2036,
   output        cfg_din2037,
   output        cfg_din2038,
   output        cfg_din2039,
   output        cfg_din2040,
   output        cfg_din2041,
   output        cfg_din2042,
   output        cfg_din2043,
   output        cfg_din2044,
   output        cfg_din2045,
   output        cfg_din2046,
   output        cfg_din2047,
   output        cfg_din2048,
   output        cfg_din2049,
   output        cfg_din2050,
   output        cfg_din2051,
   output        cfg_din2052,
   output        cfg_din2053,
   output        cfg_din2054,
   output        cfg_din2055,
   output        cfg_din2056,
   output        cfg_din2057,
   output        cfg_din2058,
   output        cfg_din2059,
   output        cfg_din2060,
   output        cfg_din2061,
   output        cfg_din2062,
   output        cfg_din2063,
   output        cfg_din2064,
   output        cfg_din2065,
   output        cfg_din2066,
   output        cfg_din2067,
   output        cfg_din2068,
   output        cfg_din2069,
   output        cfg_din2070,
   output        cfg_din2071,
   output        cfg_din2072,
   output        cfg_din2073,
   output        cfg_din2074,
   output        cfg_din2075,
   output        cfg_din2076,
   output        cfg_din2077,
   output        cfg_din2078,
   output        cfg_din2079,
   output        cfg_din2080,
   output        cfg_din2081,
   output        cfg_din2082,
   output        cfg_din2083,
   output        cfg_din2084,
   output        cfg_din2085,
   output        cfg_din2086,
   output        cfg_din2087,
   output        cfg_din2088,
   output        cfg_din2089,
   output        cfg_din2090,
   output        cfg_din2091,
   output        cfg_din2092,
   output        cfg_din2093,
   output        cfg_din2094,
   output        cfg_din2095,
   output        cfg_din2096,
   output        cfg_din2097,
   output        cfg_din2098,
   output        cfg_din2099,
   output        cfg_din2100,
   output        cfg_din2101,
   output        cfg_din2102,
   output        cfg_din2103,
   output        cfg_din2104,
   output        cfg_din2105,
   output        cfg_din2106,
   output        cfg_din2107,
   output        cfg_din2108,
   output        cfg_din2109,
   output        cfg_din2110,
   output        cfg_din2111,
   output        cfg_din2112,
   output        cfg_din2113,
   output        cfg_din2114,
   output        cfg_din2115,
   output        cfg_din2116,
   output        cfg_din2117,
   output        cfg_din2118,
   output        cfg_din2119,
   output        cfg_din2120,
   output        cfg_din2121,
   output        cfg_din2122,
   output        cfg_din2123,
   output        cfg_din2124,
   output        cfg_din2125,
   output        cfg_din2126,
   output        cfg_din2127,
   output        cfg_din2128,
   output        cfg_din2129,
   output        cfg_din2130,
   output        cfg_din2131,
   output        cfg_din2132,
   output        cfg_din2133,
   output        cfg_din2134,
   output        cfg_din2135,
   output        cfg_din2136,
   output        cfg_din2137,
   output        cfg_din2138,
   output        cfg_din2139,
   output        cfg_din2140,
   output        cfg_din2141,
   output        cfg_din2142,
   output        cfg_din2143,
   output        cfg_din2144,
   output        cfg_din2145,
   output        cfg_din2146,
   output        cfg_din2147,
   output        cfg_din2148,
   output        cfg_din2149,
   output        cfg_din2150,
   output        cfg_din2151,
   output        cfg_din2152,
   output        cfg_din2153,
   output        cfg_din2154,
   output        cfg_din2155,
   output        cfg_din2156,
   output        cfg_din2157,
   output        cfg_din2158,
   output        cfg_din2159,
   output        cfg_din2160,
   output        cfg_din2161,
   output        cfg_din2162,
   output        cfg_din2163,
   output        cfg_din2164,
   output        cfg_din2165,
   output        cfg_din2166,
   output        cfg_din2167,
   output        cfg_din2168,
   output        cfg_din2169,
   output        cfg_din2170,
   output        cfg_din2171,
   output        cfg_din2172,
   output        cfg_din2173,
   output        cfg_din2174,
   output        cfg_din2175,
   output        cfg_din2176,
   output        cfg_din2177,
   output        cfg_din2178,
   output        cfg_din2179,
   output        cfg_din2180,
   output        cfg_din2181,
   output        cfg_din2182,
   output        cfg_din2183,
   output        cfg_din2184,
   output        cfg_din2185,
   output        cfg_din2186,
   output        cfg_din2187,
   output        cfg_din2188,
   output        cfg_din2189,
   output        cfg_din2190,
   output        cfg_din2191,
   output        cfg_din2192,
   output        cfg_din2193,
   output        cfg_din2194,
   output        cfg_din2195,
   output        cfg_din2196,
   output        cfg_din2197,
   output        cfg_din2198,
   output        cfg_din2199,
   output        cfg_din2200,
   output        cfg_din2201,
   output        cfg_din2202,
   output        cfg_din2203,
   output        cfg_din2204,
   output        cfg_din2205,
   output        cfg_din2206,
   output        cfg_din2207,
   output        cfg_din2208,
   output        cfg_din2209,
   output        cfg_din2210,
   output        cfg_din2211,
   output        cfg_din2212,
   output        cfg_din2213,
   output        cfg_din2214,
   output        cfg_din2215,
   output        cfg_din2216,
   output        cfg_din2217,
   output        cfg_din2218,
   output        cfg_din2219,
   output        cfg_din2220,
   output        cfg_din2221,
   output        cfg_din2222,
   output        cfg_din2223,
   output        cfg_din2224,
   output        cfg_din2225,
   output        cfg_din2226,
   output        cfg_din2227,
   output        cfg_din2228,
   output        cfg_din2229,
   output        cfg_din2230,
   output        cfg_din2231,
   output        cfg_din2232,
   output        cfg_din2233,
   output        cfg_din2234,
   output        cfg_din2235,
   output        cfg_din2236,
   output        cfg_din2237,
   output        cfg_din2238,
   output        cfg_din2239,
   output        cfg_din2240,
   output        cfg_din2241,
   output        cfg_din2242,
   output        cfg_din2243,
   output        cfg_din2244,
   output        cfg_din2245,
   output        cfg_din2246,
   output        cfg_din2247,
   output        cfg_din2248,
   output        cfg_din2249,
   output        cfg_din2250,
   output        cfg_din2251,
   output        cfg_din2252,
   output        cfg_din2253,
   output        cfg_din2254,
   output        cfg_din2255,
   output        cfg_din2256,
   output        cfg_din2257,
   output        cfg_din2258,
   output        cfg_din2259,
   output        cfg_din2260,
   output        cfg_din2261,
   output        cfg_din2262,
   output        cfg_din2263,
   output        cfg_din2264,
   output        cfg_din2265,
   output        cfg_din2266,
   output        cfg_din2267,
   output        cfg_din2268,
   output        cfg_din2269,
   output        cfg_din2270,
   output        cfg_din2271,
   output        cfg_din2272,
   output        cfg_din2273,
   output        cfg_din2274,
   output        cfg_din2275,
   output        cfg_din2276,
   output        cfg_din2277,
   output        cfg_din2278,
   output        cfg_din2279,
   output        cfg_din2280,
   output        cfg_din2281,
   output        cfg_din2282,
   output        cfg_din2283,
   output        cfg_din2284,
   output        cfg_din2285,
   output        cfg_din2286,
   output        cfg_din2287,
   output        cfg_din2288,
   output        cfg_din2289,
   output        cfg_din2290,
   output        cfg_din2291,
   output        cfg_din2292,
   output        cfg_din2293,
   output        cfg_din2294,
   output        cfg_din2295,
   output        cfg_din2296,
   output        cfg_din2297,
   output        cfg_din2298,
   output        cfg_din2299,
   output        cfg_din2300,
   output        cfg_din2301,
   output        cfg_din2302,
   output        cfg_din2303,
   output        cfg_din2304,
   output        cfg_din2305,
   output        cfg_din2306,
   output        cfg_din2307,
   output        cfg_din2308,
   output        cfg_din2309,
   output        cfg_din2310,
   output        cfg_din2311,
   output        cfg_din2312,
   output        cfg_din2313,
   output        cfg_din2314,
   output        cfg_din2315,
   output        cfg_din2316,
   output        cfg_din2317,
   output        cfg_din2318,
   output        cfg_din2319,
   output        cfg_din2320,
   output        cfg_din2321,
   output        cfg_din2322,
   output        cfg_din2323,
   output        cfg_din2324,
   output        cfg_din2325,
   output        cfg_din2326,
   output        cfg_din2327,
   output        cfg_din2328,
   output        cfg_din2329,
   output        cfg_din2330,
   output        cfg_din2331,
   output        cfg_din2332,
   output        cfg_din2333,
   output        cfg_din2334,
   output        cfg_din2335,
   output        cfg_din2336,
   output        cfg_din2337,
   output        cfg_din2338,
   output        cfg_din2339,
   output        cfg_din2340,
   output        cfg_din2341,
   output        cfg_din2342,
   output        cfg_din2343,
   output        cfg_din2344,
   output        cfg_din2345,
   output        cfg_din2346,
   output        cfg_din2347,
   output        cfg_din2348,
   output        cfg_din2349,
   output        cfg_din2350,
   output        cfg_din2351,
   output        cfg_din2352,
   output        cfg_din2353,
   output        cfg_din2354,
   output        cfg_din2355,
   output        cfg_din2356,
   output        cfg_din2357,
   output        cfg_din2358,
   output        cfg_din2359,
   output        cfg_din2360,
   output        cfg_din2361,
   output        cfg_din2362,
   output        cfg_din2363,
   output        cfg_din2364,
   output        cfg_din2365,
   output        cfg_din2366,
   output        cfg_din2367,
   output        cfg_din2368,
   output        cfg_din2369,
   output        cfg_din2370,
   output        cfg_din2371,
   output        cfg_din2372,
   output        cfg_din2373,
   output        cfg_din2374,
   output        cfg_din2375,
   output        cfg_din2376,
   output        cfg_din2377,
   output        cfg_din2378,
   output        cfg_din2379,
   output        cfg_din2380,
   output        cfg_din2381,
   output        cfg_din2382,
   output        cfg_din2383,
   output        cfg_din2384,
   output        cfg_din2385,
   output        cfg_din2386,
   output        cfg_din2387,
   output        cfg_din2388,
   output        cfg_din2389,
   output        cfg_din2390,
   output        cfg_din2391,
   output        cfg_din2392,
   output        cfg_din2393,
   output        cfg_din2394,
   output        cfg_din2395,
   output        cfg_din2396,
   output        cfg_din2397,
   output        cfg_din2398,
   output        cfg_din2399,
   output        cfg_din2400,
   output        cfg_din2401,
   output        cfg_din2402,
   output        cfg_din2403,
   output        cfg_din2404,
   output        cfg_din2405,
   output        cfg_din2406,
   output        cfg_din2407,
   output        cfg_din2408,
   output        cfg_din2409,
   output        cfg_din2410,
   output        cfg_din2411,
   output        cfg_din2412,
   output        cfg_din2413,
   output        cfg_din2414,
   output        cfg_din2415,
   output        cfg_din2416,
   output        cfg_din2417,
   output        cfg_din2418,
   output        cfg_din2419,
   output        cfg_din2420,
   output        cfg_din2421,
   output        cfg_din2422,
   output        cfg_din2423,
   output        cfg_din2424,
   output        cfg_din2425,
   output        cfg_din2426,
   output        cfg_din2427,
   output        cfg_din2428,
   output        cfg_din2429,
   output        cfg_din2430,
   output        cfg_din2431,
   output        cfg_din2432,
   output        cfg_din2433,
   output        cfg_din2434,
   output        cfg_din2435,
   output        cfg_din2436,
   output        cfg_din2437,
   output        cfg_din2438,
   output        cfg_din2439,
   output        cfg_din2440,
   output        cfg_din2441,
   output        cfg_din2442,
   output        cfg_din2443,
   output        cfg_din2444,
   output        cfg_din2445,
   output        cfg_din2446,
   output        cfg_din2447,
   output        cfg_din2448,
   output        cfg_din2449,
   output        cfg_din2450,
   output        cfg_din2451,
   output        cfg_din2452,
   output        cfg_din2453,
   output        cfg_din2454,
   output        cfg_din2455,
   output        cfg_din2456,
   output        cfg_din2457,
   output        cfg_din2458,
   output        cfg_din2459,
   output        cfg_din2460,
   output        cfg_din2461,
   output        cfg_din2462,
   output        cfg_din2463,
   output        cfg_din2464,
   output        cfg_din2465,
   output        cfg_din2466,
   output        cfg_din2467,
   output        cfg_din2468,
   output        cfg_din2469,
   output        cfg_din2470,
   output        cfg_din2471,
   output        cfg_din2472,
   output        cfg_din2473,
   output        cfg_din2474,
   output        cfg_din2475,
   output        cfg_din2476,
   output        cfg_din2477,
   output        cfg_din2478,
   output        cfg_din2479,
   output        cfg_din2480,
   output        cfg_din2481,
   output        cfg_din2482,
   output        cfg_din2483,
   output        cfg_din2484,
   output        cfg_din2485,
   output        cfg_din2486,
   output        cfg_din2487,
   output        cfg_din2488,
   output        cfg_din2489,
   output        cfg_din2490,
   output        cfg_din2491,
   output        cfg_din2492,
   output        cfg_din2493,
   output        cfg_din2494,
   output        cfg_din2495,
   output        cfg_din2496,
   output        cfg_din2497,
   output        cfg_din2498,
   output        cfg_din2499,
   output        cfg_din2500,
   output        cfg_din2501,
   output        cfg_din2502,
   output        cfg_din2503,
   output        cfg_din2504,
   output        cfg_din2505,
   output        cfg_din2506,
   output        cfg_din2507,
   output        cfg_din2508,
   output        cfg_din2509,
   output        cfg_din2510,
   output        cfg_din2511,
   output        cfg_din2512,
   output        cfg_din2513,
   output        cfg_din2514,
   output        cfg_din2515,
   output        cfg_din2516,
   output        cfg_din2517,
   output        cfg_din2518,
   output        cfg_din2519,
   output        cfg_din2520,
   output        cfg_din2521,
   output        cfg_din2522,
   output        cfg_din2523,
   output        cfg_din2524,
   output        cfg_din2525,
   output        cfg_din2526,
   output        cfg_din2527,
   output        cfg_din2528,
   output        cfg_din2529,
   output        cfg_din2530,
   output        cfg_din2531,
   output        cfg_din2532,
   output        cfg_din2533,
   output        cfg_din2534,
   output        cfg_din2535,
   output        cfg_din2536,
   output        cfg_din2537,
   output        cfg_din2538,
   output        cfg_din2539,
   output        cfg_din2540,
   output        cfg_din2541,
   output        cfg_din2542,
   output        cfg_din2543,
   output        cfg_din2544,
   output        cfg_din2545,
   output        cfg_din2546,
   output        cfg_din2547,
   output        cfg_din2548,
   output        cfg_din2549,
   output        cfg_din2550,
   output        cfg_din2551,
   output        cfg_din2552,
   output        cfg_din2553,
   output        cfg_din2554,
   output        cfg_din2555,
   output        cfg_din2556,
   output        cfg_din2557,
   output        cfg_din2558,
   output        cfg_din2559,
   output        cfg_din2560,
   output        cfg_din2561,
   output        cfg_din2562,
   output        cfg_din2563,
   output        cfg_din2564,
   output        cfg_din2565,
   output        cfg_din2566,
   output        cfg_din2567,
   output        cfg_din2568,
   output        cfg_din2569,
   output        cfg_din2570,
   output        cfg_din2571,
   output        cfg_din2572,
   output        cfg_din2573,
   output        cfg_din2574,
   output        cfg_din2575,
   output        cfg_din2576,
   output        cfg_din2577,
   output        cfg_din2578,
   output        cfg_din2579,
   output        cfg_din2580,
   output        cfg_din2581,
   output        cfg_din2582,
   output        cfg_din2583,
   output        cfg_din2584,
   output        cfg_din2585,
   output        cfg_din2586,
   output        cfg_din2587,
   output        cfg_din2588,
   output        cfg_din2589,
   output        cfg_din2590,
   output        cfg_din2591,
   output        cfg_din2592,
   output        cfg_din2593,
   output        cfg_din2594,
   output        cfg_din2595,
   output        cfg_din2596,
   output        cfg_din2597,
   output        cfg_din2598,
   output        cfg_din2599,
   output        cfg_din2600,
   output        cfg_din2601,
   output        cfg_din2602,
   output        cfg_din2603,
   output        cfg_din2604,
   output        cfg_din2605,
   output        cfg_din2606,
   output        cfg_din2607,
   output        cfg_din2608,
   output        cfg_din2609,
   output        cfg_din2610,
   output        cfg_din2611,
   output        cfg_din2612,
   output        cfg_din2613,
   output        cfg_din2614,
   output        cfg_din2615,
   output        cfg_din2616,
   output        cfg_din2617,
   output        cfg_din2618,
   output        cfg_din2619,
   output        cfg_din2620,
   output        cfg_din2621,
   output        cfg_din2622,
   output        cfg_din2623,
   output        cfg_din2624,
   output        cfg_din2625,
   output        cfg_din2626,
   output        cfg_din2627,
   output        cfg_din2628,
   output        cfg_din2629,
   output        cfg_din2630,
   output        cfg_din2631,
   output        cfg_din2632,
   output        cfg_din2633,
   output        cfg_din2634,
   output        cfg_din2635,
   output        cfg_din2636,
   output        cfg_din2637,
   output        cfg_din2638,
   output        cfg_din2639,
   output        cfg_din2640,
   output        cfg_din2641,
   output        cfg_din2642,
   output        cfg_din2643,
   output        cfg_din2644,
   output        cfg_din2645,
   output        cfg_din2646,
   output        cfg_din2647,
   output        cfg_din2648,
   output        cfg_din2649,
   output        cfg_din2650,
   output        cfg_din2651,
   output        cfg_din2652,
   output        cfg_din2653,
   output        cfg_din2654,
   output        cfg_din2655,
   output        cfg_din2656,
   output        cfg_din2657,
   output        cfg_din2658,
   output        cfg_din2659,
   output        cfg_din2660,
   output        cfg_din2661,
   output        cfg_din2662,
   output        cfg_din2663,
   output        cfg_din2664,
   output        cfg_din2665,
   output        cfg_din2666,
   output        cfg_din2667,
   output        cfg_din2668,
   output        cfg_din2669,
   output        cfg_din2670,
   output        cfg_din2671,
   output        cfg_din2672,
   output        cfg_din2673,
   output        cfg_din2674,
   output        cfg_din2675,
   output        cfg_din2676,
   output        cfg_din2677,
   output        cfg_din2678,
   output        cfg_din2679,
   output        cfg_din2680,
   output        cfg_din2681,
   output        cfg_din2682,
   output        cfg_din2683,
   output        cfg_din2684,
   output        cfg_din2685,
   output        cfg_din2686,
   output        cfg_din2687,
   output        cfg_din2688,
   output        cfg_din2689,
   output        cfg_din2690,
   output        cfg_din2691,
   output        cfg_din2692,
   output        cfg_din2693,
   output        cfg_din2694,
   output        cfg_din2695,
   output        cfg_din2696,
   output        cfg_din2697,
   output        cfg_din2698,
   output        cfg_din2699,
   output        cfg_din2700,
   output        cfg_din2701,
   output        cfg_din2702,
   output        cfg_din2703,
   output        cfg_din2704,
   output        cfg_din2705,
   output        cfg_din2706,
   output        cfg_din2707,
   output        cfg_din2708,
   output        cfg_din2709,
   output        cfg_din2710,
   output        cfg_din2711,
   output        cfg_din2712,
   output        cfg_din2713,
   output        cfg_din2714,
   output        cfg_din2715,
   output        cfg_din2716,
   output        cfg_din2717,
   output        cfg_din2718,
   output        cfg_din2719,
   output        cfg_din2720,
   output        cfg_din2721,
   output        cfg_din2722,
   output        cfg_din2723,
   output        cfg_din2724,
   output        cfg_din2725,
   output        cfg_din2726,
   output        cfg_din2727,
   output        cfg_din2728,
   output        cfg_din2729,
   output        cfg_din2730,
   output        cfg_din2731,
   output        cfg_din2732,
   output        cfg_din2733,
   output        cfg_din2734,
   output        cfg_din2735,
   output        cfg_din2736,
   output        cfg_din2737,
   output        cfg_din2738,
   output        cfg_din2739,
   output        cfg_din2740,
   output        cfg_din2741,
   output        cfg_din2742,
   output        cfg_din2743,
   output        cfg_din2744,
   output        cfg_din2745,
   output        cfg_din2746,
   output        cfg_din2747,
   output        cfg_din2748,
   output        cfg_din2749,
   output        cfg_din2750,
   output        cfg_din2751,
   output        cfg_din2752,
   output        cfg_din2753,
   output        cfg_din2754,
   output        cfg_din2755,
   output        cfg_din2756,
   output        cfg_din2757,
   output        cfg_din2758,
   output        cfg_din2759,
   output        cfg_din2760,
   output        cfg_din2761,
   output        cfg_din2762,
   output        cfg_din2763,
   output        cfg_din2764,
   output        cfg_din2765,
   output        cfg_din2766,
   output        cfg_din2767,
   output        cfg_din2768,
   output        cfg_din2769,
   output        cfg_din2770,
   output        cfg_din2771,
   output        cfg_din2772,
   output        cfg_din2773,
   output        cfg_din2774,
   output        cfg_din2775,
   output        cfg_din2776,
   output        cfg_din2777,
   output        cfg_din2778,
   output        cfg_din2779,
   output        cfg_din2780,
   output        cfg_din2781,
   output        cfg_din2782,
   output        cfg_din2783,
   output        cfg_din2784,
   output        cfg_din2785,
   output        cfg_din2786,
   output        cfg_din2787,
   output        cfg_din2788,
   output        cfg_din2789,
   output        cfg_din2790,
   output        cfg_din2791,
   output        cfg_din2792,
   output        cfg_din2793,
   output        cfg_din2794,
   output        cfg_din2795,
   output        cfg_din2796,
   output        cfg_din2797,
   output        cfg_din2798,
   output        cfg_din2799,
   output        cfg_din2800,
   output        cfg_din2801,
   output        cfg_din2802,
   output        cfg_din2803,
   output        cfg_din2804,
   output        cfg_din2805,
   output        cfg_din2806,
   output        cfg_din2807,
   output        cfg_din2808,
   output        cfg_din2809,
   output        cfg_din2810,
   output        cfg_din2811,
   output        cfg_din2812,
   output        cfg_din2813,
   output        cfg_din2814,
   output        cfg_din2815,
   output        cfg_din2816,
   output        cfg_din2817,
   output        cfg_din2818,
   output        cfg_din2819,
   output        cfg_din2820,
   output        cfg_din2821,
   output        cfg_din2822,
   output        cfg_din2823,
   output        cfg_din2824,
   output        cfg_din2825,
   output        cfg_din2826,
   output        cfg_din2827,
   output        cfg_din2828,
   output        cfg_din2829,
   output        cfg_din2830,
   output        cfg_din2831,
   output        cfg_din2832,
   output        cfg_din2833,
   output        cfg_din2834,
   output        cfg_din2835,
   output        cfg_din2836,
   output        cfg_din2837,
   output        cfg_din2838,
   output        cfg_din2839,
   output        cfg_din2840,
   output        cfg_din2841,
   output        cfg_din2842,
   output        cfg_din2843,
   output        cfg_din2844,
   output        cfg_din2845,
   output        cfg_din2846,
   output        cfg_din2847,
   output        cfg_din2848,
   output        cfg_din2849,
   output        cfg_din2850,
   output        cfg_din2851,
   output        cfg_din2852,
   output        cfg_din2853,
   output        cfg_din2854,
   output        cfg_din2855,
   output        cfg_din2856,
   output        cfg_din2857,
   output        cfg_din2858,
   output        cfg_din2859,
   output        cfg_din2860,
   output        cfg_din2861,
   output        cfg_din2862,
   output        cfg_din2863,
   output        cfg_din2864,
   output        cfg_din2865,
   output        cfg_din2866,
   output        cfg_din2867,
   output        cfg_din2868,
   output        cfg_din2869,
   output        cfg_din2870,
   output        cfg_din2871,
   output        cfg_din2872,
   output        cfg_din2873,
   output        cfg_din2874,
   output        cfg_din2875,
   output        cfg_din2876,
   output        cfg_din2877,
   output        cfg_din2878,
   output        cfg_din2879,
   output        cfg_din2880,
   output        cfg_din2881,
   output        cfg_din2882,
   output        cfg_din2883,
   output        cfg_din2884,
   output        cfg_din2885,
   output        cfg_din2886,
   output        cfg_din2887,
   output        cfg_din2888,
   output        cfg_din2889,
   output        cfg_din2890,
   output        cfg_din2891,
   output        cfg_din2892,
   output        cfg_din2893,
   output        cfg_din2894,
   output        cfg_din2895,
   output        cfg_din2896,
   output        cfg_din2897,
   output        cfg_din2898,
   output        cfg_din2899,
   output        cfg_din2900,
   output        cfg_din2901,
   output        cfg_din2902,
   output        cfg_din2903,
   output        cfg_din2904,
   output        cfg_din2905,
   output        cfg_din2906,
   output        cfg_din2907,
   output        cfg_din2908,
   output        cfg_din2909,
   output        cfg_din2910,
   output        cfg_din2911,
   output        cfg_din2912,
   output        cfg_din2913,
   output        cfg_din2914,
   output        cfg_din2915,
   output        cfg_din2916,
   output        cfg_din2917,
   output        cfg_din2918,
   output        cfg_din2919,
   output        cfg_din2920,
   output        cfg_din2921,
   output        cfg_din2922,
   output        cfg_din2923,
   output        cfg_din2924,
   output        cfg_din2925,
   output        cfg_din2926,
   output        cfg_din2927,
   output        cfg_din2928,
   output        cfg_din2929,
   output        cfg_din2930,
   output        cfg_din2931,
   output        cfg_din2932,
   output        cfg_din2933,
   output        cfg_din2934,
   output        cfg_din2935,
   output        cfg_din2936,
   output        cfg_din2937,
   output        cfg_din2938,
   output        cfg_din2939,
   output        cfg_din2940,
   output        cfg_din2941,
   output        cfg_din2942,
   output        cfg_din2943,
   output        cfg_din2944,
   output        cfg_din2945,
   output        cfg_din2946,
   output        cfg_din2947,
   output        cfg_din2948,
   output        cfg_din2949,
   output        cfg_din2950,
   output        cfg_din2951,
   output        cfg_din2952,
   output        cfg_din2953,
   output        cfg_din2954,
   output        cfg_din2955,
   output        cfg_din2956,
   output        cfg_din2957,
   output        cfg_din2958,
   output        cfg_din2959,
   output        cfg_din2960,
   output        cfg_din2961,
   output        cfg_din2962,
   output        cfg_din2963,
   output        cfg_din2964,
   output        cfg_din2965,
   output        cfg_din2966,
   output        cfg_din2967,
   output        cfg_din2968,
   output        cfg_din2969,
   output        cfg_din2970,
   output        cfg_din2971,
   output        cfg_din2972,
   output        cfg_din2973,
   output        cfg_din2974,
   output        cfg_din2975,
   output        cfg_din2976,
   output        cfg_din2977,
   output        cfg_din2978,
   output        cfg_din2979,
   output        cfg_din2980,
   output        cfg_din2981,
   output        cfg_din2982,
   output        cfg_din2983,
   output        cfg_din2984,
   output        cfg_din2985,
   output        cfg_din2986,
   output        cfg_din2987,
   output        cfg_din2988,
   output        cfg_din2989,
   output        cfg_din2990,
   output        cfg_din2991,
   output        cfg_din2992,
   output        cfg_din2993,
   output        cfg_din2994,
   output        cfg_din2995,
   output        cfg_din2996,
   output        cfg_din2997,
   output        cfg_din2998,
   output        cfg_din2999,
   output        cfg_din3000,
   output        cfg_din3001,
   output        cfg_din3002,
   output        cfg_din3003,
   output        cfg_din3004,
   output        cfg_din3005,
   output        cfg_din3006,
   output        cfg_din3007,
   output        cfg_din3008,
   output        cfg_din3009,
   output        cfg_din3010,
   output        cfg_din3011,
   output        cfg_din3012,
   output        cfg_din3013,
   output        cfg_din3014,
   output        cfg_din3015,
   output        cfg_din3016,
   output        cfg_din3017,
   output        cfg_din3018,
   output        cfg_din3019,
   output        cfg_din3020,
   output        cfg_din3021,
   output        cfg_din3022,
   output        cfg_din3023,
   output        cfg_din3024,
   output        cfg_din3025,
   output        cfg_din3026,
   output        cfg_din3027,
   output        cfg_din3028,
   output        cfg_din3029,
   output        cfg_din3030,
   output        cfg_din3031,
   output        cfg_din3032,
   output        cfg_din3033,
   output        cfg_din3034,
   output        cfg_din3035,
   output        cfg_din3036,
   output        cfg_din3037,
   output        cfg_din3038,
   output        cfg_din3039,
   output        cfg_din3040,
   output        cfg_din3041,
   output        cfg_din3042,
   output        cfg_din3043,
   output        cfg_din3044,
   output        cfg_din3045,
   output        cfg_din3046,
   output        cfg_din3047,
   output        cfg_din3048,
   output        cfg_din3049,
   output        cfg_din3050,
   output        cfg_din3051,
   output        cfg_din3052,
   output        cfg_din3053,
   output        cfg_din3054,
   output        cfg_din3055,
   output        cfg_din3056,
   output        cfg_din3057,
   output        cfg_din3058,
   output        cfg_din3059,
   output        cfg_din3060,
   output        cfg_din3061,
   output        cfg_din3062,
   output        cfg_din3063,
   output        cfg_din3064,
   output        cfg_din3065,
   output        cfg_din3066,
   output        cfg_din3067,
   output        cfg_din3068,
   output        cfg_din3069,
   output        cfg_din3070,
   output        cfg_din3071,
   output        cfg_din3072,
   output        cfg_din3073,
   output        cfg_din3074,
   output        cfg_din3075,
   output        cfg_din3076,
   output        cfg_din3077,
   output        cfg_din3078,
   output        cfg_din3079,
   output        cfg_din3080,
   output        cfg_din3081,
   output        cfg_din3082,
   output        cfg_din3083,
   output        cfg_din3084,
   output        cfg_din3085,
   output        cfg_din3086,
   output        cfg_din3087,
   output        cfg_din3088,
   output        cfg_din3089,
   output        cfg_din3090,
   output        cfg_din3091,
   output        cfg_din3092,
   output        cfg_din3093,
   output        cfg_din3094,
   output        cfg_din3095,
   output        cfg_din3096,
   output        cfg_din3097,
   output        cfg_din3098,
   output        cfg_din3099,
   output        cfg_din3100,
   output        cfg_din3101,
   output        cfg_din3102,
   output        cfg_din3103,
   output        cfg_din3104,
   output        cfg_din3105,
   output        cfg_din3106,
   output        cfg_din3107,
   output        cfg_din3108,
   output        cfg_din3109,
   output        cfg_din3110,
   output        cfg_din3111,
   output        cfg_din3112,
   output        cfg_din3113,
   output        cfg_din3114,
   output        cfg_din3115,
   output        cfg_din3116,
   output        cfg_din3117,
   output        cfg_din3118,
   output        cfg_din3119,
   output        cfg_din3120,
   output        cfg_din3121,
   output        cfg_din3122,
   output        cfg_din3123,
   output        cfg_din3124,
   output        cfg_din3125,
   output        cfg_din3126,
   output        cfg_din3127,
   output        cfg_din3128,
   output        cfg_din3129,
   output        cfg_din3130,
   output        cfg_din3131,
   output        cfg_din3132,
   output        cfg_din3133,
   output        cfg_din3134,
   output        cfg_din3135,
   output        cfg_din3136,
   output        cfg_din3137,
   output        cfg_din3138,
   output        cfg_din3139,
   output        cfg_din3140,
   output        cfg_din3141,
   output        cfg_din3142,
   output        cfg_din3143,
   output        cfg_din3144,
   output        cfg_din3145,
   output        cfg_din3146,
   output        cfg_din3147,
   output        cfg_din3148,
   output        cfg_din3149,
   output        cfg_din3150,
   output        cfg_din3151,
   output        cfg_din3152,
   output        cfg_din3153,
   output        cfg_din3154,
   output        cfg_din3155,
   output        cfg_din3156,
   output        cfg_din3157,
   output        cfg_din3158,
   output        cfg_din3159,
   output        cfg_din3160,
   output        cfg_din3161,
   output        cfg_din3162,
   output        cfg_din3163,
   output        cfg_din3164,
   output        cfg_din3165,
   output        cfg_din3166,
   output        cfg_din3167,
   output        cfg_din3168,
   output        cfg_din3169,
   output        cfg_din3170,
   output        cfg_din3171,
   output        cfg_din3172,
   output        cfg_din3173,
   output        cfg_din3174,
   output        cfg_din3175,
   output        cfg_din3176,
   output        cfg_din3177,
   output        cfg_din3178,
   output        cfg_din3179,
   output        cfg_din3180,
   output        cfg_din3181,
   output        cfg_din3182,
   output        cfg_din3183,
   output        cfg_din3184,
   output        cfg_din3185,
   output        cfg_din3186,
   output        cfg_din3187,
   output        cfg_din3188,
   output        cfg_din3189,
   output        cfg_din3190,
   output        cfg_din3191,
   output        cfg_din3192,
   output        cfg_din3193,
   output        cfg_din3194,
   output        cfg_din3195,
   output        cfg_din3196,
   output        cfg_din3197,
   output        cfg_din3198,
   output        cfg_din3199,
   output        cfg_din3200,
   output        cfg_din3201,
   output        cfg_din3202,
   output        cfg_din3203,
   output        cfg_din3204,
   output        cfg_din3205,
   output        cfg_din3206,
   output        cfg_din3207,
   output        cfg_din3208,
   output        cfg_din3209,
   output        cfg_din3210,
   output        cfg_din3211,
   output        cfg_din3212,
   output        cfg_din3213,
   output        cfg_din3214,
   output        cfg_din3215,
   output        cfg_din3216,
   output        cfg_din3217,
   output        cfg_din3218,
   output        cfg_din3219,
   output        cfg_din3220,
   output        cfg_din3221,
   output        cfg_din3222,
   output        cfg_din3223,
   output        cfg_din3224,
   output        cfg_din3225,
   output        cfg_din3226,
   output        cfg_din3227,
   output        cfg_din3228,
   output        cfg_din3229,
   output        cfg_din3230,
   output        cfg_din3231,
   output        cfg_din3232,
   output        cfg_din3233,
   output        cfg_din3234,
   output        cfg_din3235,
   output        cfg_din3236,
   output        cfg_din3237,
   output        cfg_din3238,
   output        cfg_din3239,
   output        cfg_din3240,
   output        cfg_din3241,
   output        cfg_din3242,
   output        cfg_din3243,
   output        cfg_din3244,
   output        cfg_din3245,
   output        cfg_din3246,
   output        cfg_din3247,
   output        cfg_din3248,
   output        cfg_din3249,
   output        cfg_din3250,
   output        cfg_din3251,
   output        cfg_din3252,
   output        cfg_din3253,
   output        cfg_din3254,
   output        cfg_din3255,
   output        cfg_din3256,
   output        cfg_din3257,
   output        cfg_din3258,
   output        cfg_din3259,
   output        cfg_din3260,
   output        cfg_din3261,
   output        cfg_din3262,
   output        cfg_din3263,
   output        cfg_din3264,
   output        cfg_din3265,
   output        cfg_din3266,
   output        cfg_din3267,
   output        cfg_din3268,
   output        cfg_din3269,
   output        cfg_din3270,
   output        cfg_din3271,
   output        cfg_din3272,
   output        cfg_din3273,
   output        cfg_din3274,
   output        cfg_din3275,
   output        cfg_din3276,
   output        cfg_din3277,
   output        cfg_din3278,
   output        cfg_din3279,
   output        cfg_din3280,
   output        cfg_din3281,
   output        cfg_din3282,
   output        cfg_din3283,
   output        cfg_din3284,
   output        cfg_din3285,
   output        cfg_din3286,
   output        cfg_din3287,
   output        cfg_din3288,
   output        cfg_din3289,
   output        cfg_din3290,
   output        cfg_din3291,
   output        cfg_din3292,
   output        cfg_din3293,
   output        cfg_din3294,
   output        cfg_din3295,
   output        cfg_din3296,
   output        cfg_din3297,
   output        cfg_din3298,
   output        cfg_din3299,
   output        cfg_din3300,
   output        cfg_din3301,
   output        cfg_din3302,
   output        cfg_din3303,
   output        cfg_din3304,
   output        cfg_din3305,
   output        cfg_din3306,
   output        cfg_din3307,
   output        cfg_din3308,
   output        cfg_din3309,
   output        cfg_din3310,
   output        cfg_din3311,
   output        cfg_din3312,
   output        cfg_din3313,
   output        cfg_din3314,
   output        cfg_din3315,
   output        cfg_din3316,
   output        cfg_din3317,
   output        cfg_din3318,
   output        cfg_din3319,
   output        cfg_din3320,
   output        cfg_din3321,
   output        cfg_din3322,
   output        cfg_din3323,
   output        cfg_din3324,
   output        cfg_din3325,
   output        cfg_din3326,
   output        cfg_din3327,
   output        cfg_din3328,
   output        cfg_din3329,
   output        cfg_din3330,
   output        cfg_din3331,
   output        cfg_din3332,
   output        cfg_din3333,
   output        cfg_din3334,
   output        cfg_din3335,
   output        cfg_din3336,
   output        cfg_din3337,
   output        cfg_din3338,
   output        cfg_din3339,
   output        cfg_din3340,
   output        cfg_din3341,
   output        cfg_din3342,
   output        cfg_din3343,
   output        cfg_din3344,
   output        cfg_din3345,
   output        cfg_din3346,
   output        cfg_din3347,
   output        cfg_din3348,
   output        cfg_din3349,
   output        cfg_din3350,
   output        cfg_din3351,
   output        cfg_din3352,
   output        cfg_din3353,
   output        cfg_din3354,
   output        cfg_din3355,
   output        cfg_din3356,
   output        cfg_din3357,
   output        cfg_din3358,
   output        cfg_din3359,
   output        cfg_din3360,
   output        cfg_din3361,
   output        cfg_din3362,
   output        cfg_din3363,
   output        cfg_din3364,
   output        cfg_din3365,
   output        cfg_din3366,
   output        cfg_din3367,
   output        cfg_din3368,
   output        cfg_din3369,
   output        cfg_din3370,
   output        cfg_din3371,
   output        cfg_din3372,
   output        cfg_din3373,
   output        cfg_din3374,
   output        cfg_din3375,
   output        cfg_din3376,
   output        cfg_din3377,
   output        cfg_din3378,
   output        cfg_din3379,
   output        cfg_din3380,
   output        cfg_din3381,
   output        cfg_din3382,
   output        cfg_din3383,
   output        cfg_din3384,
   output        cfg_din3385,
   output        cfg_din3386,
   output        cfg_din3387,
   output        cfg_din3388,
   output        cfg_din3389,
   output        cfg_din3390,
   output        cfg_din3391,
   output        cfg_din3392,
   output        cfg_din3393,
   output        cfg_din3394,
   output        cfg_din3395,
   output        cfg_din3396,
   output        cfg_din3397,
   output        cfg_din3398,
   output        cfg_din3399,
   output        cfg_din3400,
   output        cfg_din3401,
   output        cfg_din3402,
   output        cfg_din3403,
   output        cfg_din3404,
   output        cfg_din3405,
   output        cfg_din3406,
   output        cfg_din3407,
   output        cfg_din3408,
   output        cfg_din3409,
   output        cfg_din3410,
   output        cfg_din3411,
   output        cfg_din3412,
   output        cfg_din3413,
   output        cfg_din3414,
   output        cfg_din3415,
   output        cfg_din3416,
   output        cfg_din3417,
   output        cfg_din3418,
   output        cfg_din3419,
   output        cfg_din3420,
   output        cfg_din3421,
   output        cfg_din3422,
   output        cfg_din3423,
   output        cfg_din3424,
   output        cfg_din3425,
   output        cfg_din3426,
   output        cfg_din3427,
   output        cfg_din3428,
   output        cfg_din3429,
   output        cfg_din3430,
   output        cfg_din3431,
   output        cfg_din3432,
   output        cfg_din3433,
   output        cfg_din3434,
   output        cfg_din3435,
   output        cfg_din3436,
   output        cfg_din3437,
   output        cfg_din3438,
   output        cfg_din3439,
   output        cfg_din3440,
   output        cfg_din3441,
   output        cfg_din3442,
   output        cfg_din3443,
   output        cfg_din3444,
   output        cfg_din3445,
   output        cfg_din3446,
   output        cfg_din3447,
   output        cfg_din3448,
   output        cfg_din3449,
   output        cfg_din3450,
   output        cfg_din3451,
   output        cfg_din3452,
   output        cfg_din3453,
   output        cfg_din3454,
   output        cfg_din3455,
   output        cfg_din3456,
   output        cfg_din3457,
   output        cfg_din3458,
   output        cfg_din3459,
   output        cfg_din3460,
   output        cfg_din3461,
   output        cfg_din3462,
   output        cfg_din3463,
   output        cfg_din3464,
   output        cfg_din3465,
   output        cfg_din3466,
   output        cfg_din3467,
   output        cfg_din3468,
   output        cfg_din3469,
   output        cfg_din3470,
   output        cfg_din3471,
   output        cfg_din3472,
   output        cfg_din3473,
   output        cfg_din3474,
   output        cfg_din3475,
   output        cfg_din3476,
   output        cfg_din3477,
   output        cfg_din3478,
   output        cfg_din3479,
   output        cfg_din3480,
   output        cfg_din3481,
   output        cfg_din3482,
   output        cfg_din3483,
   output        cfg_din3484,
   output        cfg_din3485,
   output        cfg_din3486,
   output        cfg_din3487,
   output        cfg_din3488,
   output        cfg_din3489,
   output        cfg_din3490,
   output        cfg_din3491,
   output        cfg_din3492,
   output        cfg_din3493,
   output        cfg_din3494,
   output        cfg_din3495,
   output        cfg_din3496,
   output        cfg_din3497,
   output        cfg_din3498,
   output        cfg_din3499,
   output        cfg_din3500,
   output        cfg_din3501,
   output        cfg_din3502,
   output        cfg_din3503,
   output        cfg_din3504,
   output        cfg_din3505,
   output        cfg_din3506,
   output        cfg_din3507,
   output        cfg_din3508,
   output        cfg_din3509,
   output        cfg_din3510,
   output        cfg_din3511,
   output        cfg_din3512,
   output        cfg_din3513,
   output        cfg_din3514,
   output        cfg_din3515,
   output        cfg_din3516,
   output        cfg_din3517,
   output        cfg_din3518,
   output        cfg_din3519,
   output        cfg_din3520,
   output        cfg_din3521,
   output        cfg_din3522,
   output        cfg_din3523,
   output        cfg_din3524,
   output        cfg_din3525,
   output        cfg_din3526,
   output        cfg_din3527,
   output        cfg_din3528,
   output        cfg_din3529,
   output        cfg_din3530,
   output        cfg_din3531,
   output        cfg_din3532,
   output        cfg_din3533,
   output        cfg_din3534,
   output        cfg_din3535,
   output        cfg_din3536,
   output        cfg_din3537,
   output        cfg_din3538,
   output        cfg_din3539,
   output        cfg_din3540,
   output        cfg_din3541,
   output        cfg_din3542,
   output        cfg_din3543,
   output        cfg_din3544,
   output        cfg_din3545,
   output        cfg_din3546,
   output        cfg_din3547,
   output        cfg_din3548,
   output        cfg_din3549,
   output        cfg_din3550,
   output        cfg_din3551,
   output        cfg_din3552,
   output        cfg_din3553,
   output        cfg_din3554,
   output        cfg_din3555,
   output        cfg_din3556,
   output        cfg_din3557,
   output        cfg_din3558,
   output        cfg_din3559,
   output        cfg_din3560,
   output        cfg_din3561,
   output        cfg_din3562,
   output        cfg_din3563,
   output        cfg_din3564,
   output        cfg_din3565,
   output        cfg_din3566,
   output        cfg_din3567,
   output        cfg_din3568,
   output        cfg_din3569,
   output        cfg_din3570,
   output        cfg_din3571,
   output        cfg_din3572,
   output        cfg_din3573,
   output        cfg_din3574,
   output        cfg_din3575,
   output        cfg_din3576,
   output        cfg_din3577,
   output        cfg_din3578,
   output        cfg_din3579,
   output        cfg_din3580,
   output        cfg_din3581,
   output        cfg_din3582,
   output        cfg_din3583,
   output        cfg_din3584,
   output        cfg_din3585,
   output        cfg_din3586,
   output        cfg_din3587,
   output        cfg_din3588,
   output        cfg_din3589,
   output        cfg_din3590,
   output        cfg_din3591,
   output        cfg_din3592,
   output        cfg_din3593,
   output        cfg_din3594,
   output        cfg_din3595,
   output        cfg_din3596,
   output        cfg_din3597,
   output        cfg_din3598,
   output        cfg_din3599,
   output        cfg_din3600,
   output        cfg_din3601,
   output        cfg_din3602,
   output        cfg_din3603,
   output        cfg_din3604,
   output        cfg_din3605,
   output        cfg_din3606,
   output        cfg_din3607,
   output        cfg_din3608,
   output        cfg_din3609,
   output        cfg_din3610,
   output        cfg_din3611,
   output        cfg_din3612,
   output        cfg_din3613,
   output        cfg_din3614,
   output        cfg_din3615,
   output        cfg_din3616,
   output        cfg_din3617,
   output        cfg_din3618,
   output        cfg_din3619,
   output        cfg_din3620,
   output        cfg_din3621,
   output        cfg_din3622,
   output        cfg_din3623,
   output        cfg_din3624,
   output        cfg_din3625,
   output        cfg_din3626,
   output        cfg_din3627,
   output        cfg_din3628,
   output        cfg_din3629,
   output        cfg_din3630,
   output        cfg_din3631,
   output        cfg_din3632,
   output        cfg_din3633,
   output        cfg_din3634,
   output        cfg_din3635,
   output        cfg_din3636,
   output        cfg_din3637,
   output        cfg_din3638,
   output        cfg_din3639,
   output        cfg_din3640,
   output        cfg_din3641,
   output        cfg_din3642,
   output        cfg_din3643,
   output        cfg_din3644,
   output        cfg_din3645,
   output        cfg_din3646,
   output        cfg_din3647,
   output        cfg_din3648,
   output        cfg_din3649,
   output        cfg_din3650,
   output        cfg_din3651,
   output        cfg_din3652,
   output        cfg_din3653,
   output        cfg_din3654,
   output        cfg_din3655,
   output        cfg_din3656,
   output        cfg_din3657,
   output        cfg_din3658,
   output        cfg_din3659,
   output        cfg_din3660,
   output        cfg_din3661,
   output        cfg_din3662,
   output        cfg_din3663,
   output        cfg_din3664,
   output        cfg_din3665,
   output        cfg_din3666,
   output        cfg_din3667,
   output        cfg_din3668,
   output        cfg_din3669,
   output        cfg_din3670,
   output        cfg_din3671,
   output        cfg_din3672,
   output        cfg_din3673,
   output        cfg_din3674,
   output        cfg_din3675,
   output        cfg_din3676,
   output        cfg_din3677,
   output        cfg_din3678,
   output        cfg_din3679,
   output        cfg_din3680,
   output        cfg_din3681,
   output        cfg_din3682,
   output        cfg_din3683,
   output        cfg_din3684,
   output        cfg_din3685,
   output        cfg_din3686,
   output        cfg_din3687,
   output        cfg_din3688,
   output        cfg_din3689,
   output        cfg_din3690,
   output        cfg_din3691,
   output        cfg_din3692,
   output        cfg_din3693,
   output        cfg_din3694,
   output        cfg_din3695,
   output        cfg_din3696,
   output        cfg_din3697,
   output        cfg_din3698,
   output        cfg_din3699,
   output        cfg_din3700,
   output        cfg_din3701,
   output        cfg_din3702,
   output        cfg_din3703,
   output        cfg_din3704,
   output        cfg_din3705,
   output        cfg_din3706,
   output        cfg_din3707,
   output        cfg_din3708,
   output        cfg_din3709,
   output        cfg_din3710,
   output        cfg_din3711,
   output        cfg_din3712,
   output        cfg_din3713,
   output        cfg_din3714,
   output        cfg_din3715,
   output        cfg_din3716,
   output        cfg_din3717,
   output        cfg_din3718,
   output        cfg_din3719,
   output        cfg_din3720,
   output        cfg_din3721,
   output        cfg_din3722,
   output        cfg_din3723,
   output        cfg_din3724,
   output        cfg_din3725,
   output        cfg_din3726,
   output        cfg_din3727,
   output        cfg_din3728,
   output        cfg_din3729,
   output        cfg_din3730,
   output        cfg_din3731,
   output        cfg_din3732,
   output        cfg_din3733,
   output        cfg_din3734,
   output        cfg_din3735,
   output        cfg_din3736,
   output        cfg_din3737,
   output        cfg_din3738,
   output        cfg_din3739,
   output        cfg_din3740,
   output        cfg_din3741,
   output        cfg_din3742,
   output        cfg_din3743,
   output        cfg_din3744,
   output        cfg_din3745,
   output        cfg_din3746,
   output        cfg_din3747,
   output        cfg_din3748,
   output        cfg_din3749,
   output        cfg_din3750,
   output        cfg_din3751,
   output        cfg_din3752,
   output        cfg_din3753,
   output        cfg_din3754,
   output        cfg_din3755,
   output        cfg_din3756,
   output        cfg_din3757,
   output        cfg_din3758,
   output        cfg_din3759,
   output        cfg_din3760,
   output        cfg_din3761,
   output        cfg_din3762,
   output        cfg_din3763,
   output        cfg_din3764,
   output        cfg_din3765,
   output        cfg_din3766,
   output        cfg_din3767,
   output        cfg_din3768,
   output        cfg_din3769,
   output        cfg_din3770,
   output        cfg_din3771,
   output        cfg_din3772,
   output        cfg_din3773,
   output        cfg_din3774,
   output        cfg_din3775,
   output        cfg_din3776,
   output        cfg_din3777,
   output        cfg_din3778,
   output        cfg_din3779,
   output        cfg_din3780,
   output        cfg_din3781,
   output        cfg_din3782,
   output        cfg_din3783,
   output        cfg_din3784,
   output        cfg_din3785,
   output        cfg_din3786,
   output        cfg_din3787,
   output        cfg_din3788,
   output        cfg_din3789,
   output        cfg_din3790,
   output        cfg_din3791,
   output        cfg_din3792,
   output        cfg_din3793,
   output        cfg_din3794,
   output        cfg_din3795,
   output        cfg_din3796,
   output        cfg_din3797,
   output        cfg_din3798,
   output        cfg_din3799,
   output        cfg_din3800,
   output        cfg_din3801,
   output        cfg_din3802,
   output        cfg_din3803,
   output        cfg_din3804,
   output        cfg_din3805,
   output        cfg_din3806,
   output        cfg_din3807,
   output        cfg_din3808,
   output        cfg_din3809,
   output        cfg_din3810,
   output        cfg_din3811,
   output        cfg_din3812,
   output        cfg_din3813,
   output        cfg_din3814,
   output        cfg_din3815,
   output        cfg_din3816,
   output        cfg_din3817,
   output        cfg_din3818,
   output        cfg_din3819,
   output        cfg_din3820,
   output        cfg_din3821,
   output        cfg_din3822,
   output        cfg_din3823,
   output        cfg_din3824,
   output        cfg_din3825,
   output        cfg_din3826,
   output        cfg_din3827,
   output        cfg_din3828,
   output        cfg_din3829,
   output        cfg_din3830,
   output        cfg_din3831,
   output        cfg_din3832,
   output        cfg_din3833,
   output        cfg_din3834,
   output        cfg_din3835,
   output        cfg_din3836,
   output        cfg_din3837,
   output        cfg_din3838,
   output        cfg_din3839,
   output        cfg_din3840,
   output        cfg_din3841,
   output        cfg_din3842,
   output        cfg_din3843,
   output        cfg_din3844,
   output        cfg_din3845,
   output        cfg_din3846,
   output        cfg_din3847,
   output        cfg_din3848,
   output        cfg_din3849,
   output        cfg_din3850,
   output        cfg_din3851,
   output        cfg_din3852,
   output        cfg_din3853,
   output        cfg_din3854,
   output        cfg_din3855,
   output        cfg_din3856,
   output        cfg_din3857,
   output        cfg_din3858,
   output        cfg_din3859,
   output        cfg_din3860,
   output        cfg_din3861,
   output        cfg_din3862,
   output        cfg_din3863,
   output        cfg_din3864,
   output        cfg_din3865,
   output        cfg_din3866,
   output        cfg_din3867,
   output        cfg_din3868,
   output        cfg_din3869,
   output        cfg_din3870,
   output        cfg_din3871,
   output        cfg_din3872,
   output        cfg_din3873,
   output        cfg_din3874,
   output        cfg_din3875,
   output        cfg_din3876,
   output        cfg_din3877,
   output        cfg_din3878,
   output        cfg_din3879,
   output        cfg_din3880,
   output        cfg_din3881,
   output        cfg_din3882,
   output        cfg_din3883,
   output        cfg_din3884,
   output        cfg_din3885,
   output        cfg_din3886,
   output        cfg_din3887,
   output        cfg_din3888,
   output        cfg_din3889,
   output        cfg_din3890,
   output        cfg_din3891,
   output        cfg_din3892,
   output        cfg_din3893,
   output        cfg_din3894,
   output        cfg_din3895,
   output        cfg_din3896,
   output        cfg_din3897,
   output        cfg_din3898,
   output        cfg_din3899,
   output        cfg_din3900,
   output        cfg_din3901,
   output        cfg_din3902,
   output        cfg_din3903,
   output        cfg_din3904,
   output        cfg_din3905,
   output        cfg_din3906,
   output        cfg_din3907,
   output        cfg_din3908,
   output        cfg_din3909,
   output        cfg_din3910,
   output        cfg_din3911,
   output        cfg_din3912,
   output        cfg_din3913,
   output        cfg_din3914,
   output        cfg_din3915,
   output        cfg_din3916,
   output        cfg_din3917,
   output        cfg_din3918,
   output        cfg_din3919,
   output        cfg_din3920,
   output        cfg_din3921,
   output        cfg_din3922,
   output        cfg_din3923,
   output        cfg_din3924,
   output        cfg_din3925,
   output        cfg_din3926,
   output        cfg_din3927,
   output        cfg_din3928,
   output        cfg_din3929,
   output        cfg_din3930,
   output        cfg_din3931,
   output        cfg_din3932,
   output        cfg_din3933,
   output        cfg_din3934,
   output        cfg_din3935,
   output        cfg_din3936,
   output        cfg_din3937,
   output        cfg_din3938,
   output        cfg_din3939,
   output        cfg_din3940,
   output        cfg_din3941,
   output        cfg_din3942,
   output        cfg_din3943,
   output        cfg_din3944,
   output        cfg_din3945,
   output        cfg_din3946,
   output        cfg_din3947,
   output        cfg_din3948,
   output        cfg_din3949,
   output        cfg_din3950,
   output        cfg_din3951,
   output        cfg_din3952,
   output        cfg_din3953,
   output        cfg_din3954,
   output        cfg_din3955,
   output        cfg_din3956,
   output        cfg_din3957,
   output        cfg_din3958,
   output        cfg_din3959,
   output        cfg_din3960,
   output        cfg_din3961,
   output        cfg_din3962,
   output        cfg_din3963,
   output        cfg_din3964,
   output        cfg_din3965,
   output        cfg_din3966,
   output        cfg_din3967,
   output        cfg_din3968,
   output        cfg_din3969,
   output        cfg_din3970,
   output        cfg_din3971,
   output        cfg_din3972,
   output        cfg_din3973,
   output        cfg_din3974,
   output        cfg_din3975,
   output        cfg_din3976,
   output        cfg_din3977,
   output        cfg_din3978,
   output        cfg_din3979,
   output        cfg_din3980,
   output        cfg_din3981,
   output        cfg_din3982,
   output        cfg_din3983,
   output        cfg_din3984,
   output        cfg_din3985,
   output        cfg_din3986,
   output        cfg_din3987,
   output        cfg_din3988,
   output        cfg_din3989,
   output        cfg_din3990,
   output        cfg_din3991,
   output        cfg_din3992,
   output        cfg_din3993,
   output        cfg_din3994,
   output        cfg_din3995,
   output        cfg_din3996,
   output        cfg_din3997,
   output        cfg_din3998,
   output        cfg_din3999,
   output        cfg_din4000,
   output        cfg_din4001,
   output        cfg_din4002,
   output        cfg_din4003,
   output        cfg_din4004,
   output        cfg_din4005,
   output        cfg_din4006,
   output        cfg_din4007,
   output        cfg_din4008,
   output        cfg_din4009,
   output        cfg_din4010,
   output        cfg_din4011,
   output        cfg_din4012,
   output        cfg_din4013,
   output        cfg_din4014,
   output        cfg_din4015,
   output        cfg_din4016,
   output        cfg_din4017,
   output        cfg_din4018,
   output        cfg_din4019,
   output        cfg_din4020,
   output        cfg_din4021,
   output        cfg_din4022,
   output        cfg_din4023,
   output        cfg_din4024,
   output        cfg_din4025,
   output        cfg_din4026,
   output        cfg_din4027,
   output        cfg_din4028,
   output        cfg_din4029,
   output        cfg_din4030,
   output        cfg_din4031,
   output        cfg_din4032,
   output        cfg_din4033,
   output        cfg_din4034,
   output        cfg_din4035,
   output        cfg_din4036,
   output        cfg_din4037,
   output        cfg_din4038,
   output        cfg_din4039,
   output        cfg_din4040,
   output        cfg_din4041,
   output        cfg_din4042,
   output        cfg_din4043,
   output        cfg_din4044,
   output        cfg_din4045,
   output        cfg_din4046,
   output        cfg_din4047,
   output        cfg_din4048,
   output        cfg_din4049,
   output        cfg_din4050,
   output        cfg_din4051,
   output        cfg_din4052,
   output        cfg_din4053,
   output        cfg_din4054,
   output        cfg_din4055,
   output        cfg_din4056,
   output        cfg_din4057,
   output        cfg_din4058,
   output        cfg_din4059,
   output        cfg_din4060,
   output        cfg_din4061,
   output        cfg_din4062,
   output        cfg_din4063,
   output        cfg_din4064,
   output        cfg_din4065,
   output        cfg_din4066,
   output        cfg_din4067,
   output        cfg_din4068,
   output        cfg_din4069,
   output        cfg_din4070,
   output        cfg_din4071,
   output        cfg_din4072,
   output        cfg_din4073,
   output        cfg_din4074,
   output        cfg_din4075,
   output        cfg_din4076,
   output        cfg_din4077,
   output        cfg_din4078,
   output        cfg_din4079,
   output        cfg_din4080,
   output        cfg_din4081,
   output        cfg_din4082,
   output        cfg_din4083,
   output        cfg_din4084,
   output        cfg_din4085,
   output        cfg_din4086,
   output        cfg_din4087,
   output        cfg_din4088,
   output        cfg_din4089,
   output        cfg_din4090,
   output        cfg_din4091,
   output        cfg_din4092,
   output        cfg_din4093,
   output        cfg_din4094,
   output        cfg_din4095,
   output        tc_cfg_din,
   output        cc_cfg_din0,
   output        cc_cfg_din1,
   output        cc_cfg_din2,
   output        cc_cfg_din3,

